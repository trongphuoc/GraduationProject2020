// soc_system.v

// Generated using ACDS version 13.0sp1 232 at 2013.08.29.23:21:29

`timescale 1 ps / 1 ps
module soc_system (
		input  wire        reset_reset_n,                             //                          reset.reset_n
		output wire [14:0] memory_mem_a,                              //                         memory.mem_a
		output wire [2:0]  memory_mem_ba,                             //                               .mem_ba
		output wire        memory_mem_ck,                             //                               .mem_ck
		output wire        memory_mem_ck_n,                           //                               .mem_ck_n
		output wire        memory_mem_cke,                            //                               .mem_cke
		output wire        memory_mem_cs_n,                           //                               .mem_cs_n
		output wire        memory_mem_ras_n,                          //                               .mem_ras_n
		output wire        memory_mem_cas_n,                          //                               .mem_cas_n
		output wire        memory_mem_we_n,                           //                               .mem_we_n
		output wire        memory_mem_reset_n,                        //                               .mem_reset_n
		inout  wire [31:0] memory_mem_dq,                             //                               .mem_dq
		inout  wire [3:0]  memory_mem_dqs,                            //                               .mem_dqs
		inout  wire [3:0]  memory_mem_dqs_n,                          //                               .mem_dqs_n
		output wire        memory_mem_odt,                            //                               .mem_odt
		output wire [3:0]  memory_mem_dm,                             //                               .mem_dm
		input  wire        memory_oct_rzqin,                          //                               .oct_rzqin
		output wire        hps_0_hps_io_hps_io_emac1_inst_TX_CLK,     //                   hps_0_hps_io.hps_io_emac1_inst_TX_CLK
		output wire        hps_0_hps_io_hps_io_emac1_inst_TXD0,       //                               .hps_io_emac1_inst_TXD0
		output wire        hps_0_hps_io_hps_io_emac1_inst_TXD1,       //                               .hps_io_emac1_inst_TXD1
		output wire        hps_0_hps_io_hps_io_emac1_inst_TXD2,       //                               .hps_io_emac1_inst_TXD2
		output wire        hps_0_hps_io_hps_io_emac1_inst_TXD3,       //                               .hps_io_emac1_inst_TXD3
		input  wire        hps_0_hps_io_hps_io_emac1_inst_RXD0,       //                               .hps_io_emac1_inst_RXD0
		inout  wire        hps_0_hps_io_hps_io_emac1_inst_MDIO,       //                               .hps_io_emac1_inst_MDIO
		output wire        hps_0_hps_io_hps_io_emac1_inst_MDC,        //                               .hps_io_emac1_inst_MDC
		input  wire        hps_0_hps_io_hps_io_emac1_inst_RX_CTL,     //                               .hps_io_emac1_inst_RX_CTL
		output wire        hps_0_hps_io_hps_io_emac1_inst_TX_CTL,     //                               .hps_io_emac1_inst_TX_CTL
		input  wire        hps_0_hps_io_hps_io_emac1_inst_RX_CLK,     //                               .hps_io_emac1_inst_RX_CLK
		input  wire        hps_0_hps_io_hps_io_emac1_inst_RXD1,       //                               .hps_io_emac1_inst_RXD1
		input  wire        hps_0_hps_io_hps_io_emac1_inst_RXD2,       //                               .hps_io_emac1_inst_RXD2
		input  wire        hps_0_hps_io_hps_io_emac1_inst_RXD3,       //                               .hps_io_emac1_inst_RXD3
		inout  wire        hps_0_hps_io_hps_io_qspi_inst_IO0,         //                               .hps_io_qspi_inst_IO0
		inout  wire        hps_0_hps_io_hps_io_qspi_inst_IO1,         //                               .hps_io_qspi_inst_IO1
		inout  wire        hps_0_hps_io_hps_io_qspi_inst_IO2,         //                               .hps_io_qspi_inst_IO2
		inout  wire        hps_0_hps_io_hps_io_qspi_inst_IO3,         //                               .hps_io_qspi_inst_IO3
		output wire        hps_0_hps_io_hps_io_qspi_inst_SS0,         //                               .hps_io_qspi_inst_SS0
		output wire        hps_0_hps_io_hps_io_qspi_inst_CLK,         //                               .hps_io_qspi_inst_CLK
		inout  wire        hps_0_hps_io_hps_io_sdio_inst_CMD,         //                               .hps_io_sdio_inst_CMD
		inout  wire        hps_0_hps_io_hps_io_sdio_inst_D0,          //                               .hps_io_sdio_inst_D0
		inout  wire        hps_0_hps_io_hps_io_sdio_inst_D1,          //                               .hps_io_sdio_inst_D1
		output wire        hps_0_hps_io_hps_io_sdio_inst_CLK,         //                               .hps_io_sdio_inst_CLK
		inout  wire        hps_0_hps_io_hps_io_sdio_inst_D2,          //                               .hps_io_sdio_inst_D2
		inout  wire        hps_0_hps_io_hps_io_sdio_inst_D3,          //                               .hps_io_sdio_inst_D3
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D0,          //                               .hps_io_usb1_inst_D0
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D1,          //                               .hps_io_usb1_inst_D1
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D2,          //                               .hps_io_usb1_inst_D2
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D3,          //                               .hps_io_usb1_inst_D3
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D4,          //                               .hps_io_usb1_inst_D4
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D5,          //                               .hps_io_usb1_inst_D5
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D6,          //                               .hps_io_usb1_inst_D6
		inout  wire        hps_0_hps_io_hps_io_usb1_inst_D7,          //                               .hps_io_usb1_inst_D7
		input  wire        hps_0_hps_io_hps_io_usb1_inst_CLK,         //                               .hps_io_usb1_inst_CLK
		output wire        hps_0_hps_io_hps_io_usb1_inst_STP,         //                               .hps_io_usb1_inst_STP
		input  wire        hps_0_hps_io_hps_io_usb1_inst_DIR,         //                               .hps_io_usb1_inst_DIR
		input  wire        hps_0_hps_io_hps_io_usb1_inst_NXT,         //                               .hps_io_usb1_inst_NXT
		output wire        hps_0_hps_io_hps_io_spim1_inst_CLK,        //                               .hps_io_spim1_inst_CLK
		output wire        hps_0_hps_io_hps_io_spim1_inst_MOSI,       //                               .hps_io_spim1_inst_MOSI
		input  wire        hps_0_hps_io_hps_io_spim1_inst_MISO,       //                               .hps_io_spim1_inst_MISO
		output wire        hps_0_hps_io_hps_io_spim1_inst_SS0,        //                               .hps_io_spim1_inst_SS0
		input  wire        hps_0_hps_io_hps_io_uart0_inst_RX,         //                               .hps_io_uart0_inst_RX
		output wire        hps_0_hps_io_hps_io_uart0_inst_TX,         //                               .hps_io_uart0_inst_TX
		inout  wire        hps_0_hps_io_hps_io_i2c0_inst_SDA,         //                               .hps_io_i2c0_inst_SDA
		inout  wire        hps_0_hps_io_hps_io_i2c0_inst_SCL,         //                               .hps_io_i2c0_inst_SCL
		inout  wire        hps_0_hps_io_hps_io_i2c1_inst_SDA,         //                               .hps_io_i2c1_inst_SDA
		inout  wire        hps_0_hps_io_hps_io_i2c1_inst_SCL,         //                               .hps_io_i2c1_inst_SCL
		inout  wire        hps_0_hps_io_hps_io_gpio_inst_GPIO09,      //                               .hps_io_gpio_inst_GPIO09
		inout  wire        hps_0_hps_io_hps_io_gpio_inst_GPIO35,      //                               .hps_io_gpio_inst_GPIO35
		inout  wire        hps_0_hps_io_hps_io_gpio_inst_GPIO40,      //                               .hps_io_gpio_inst_GPIO40
		inout  wire        hps_0_hps_io_hps_io_gpio_inst_GPIO41,      //                               .hps_io_gpio_inst_GPIO41
		inout  wire        hps_0_hps_io_hps_io_gpio_inst_GPIO48,      //                               .hps_io_gpio_inst_GPIO48
		inout  wire        hps_0_hps_io_hps_io_gpio_inst_GPIO53,      //                               .hps_io_gpio_inst_GPIO53
		inout  wire        hps_0_hps_io_hps_io_gpio_inst_GPIO54,      //                               .hps_io_gpio_inst_GPIO54
		inout  wire        hps_0_hps_io_hps_io_gpio_inst_GPIO61,      //                               .hps_io_gpio_inst_GPIO61
		output wire [9:0]  led_pio_external_connection_export,        //    led_pio_external_connection.export
		input  wire [3:0]  dipsw_pio_external_connection_export,      //  dipsw_pio_external_connection.export
		input  wire [1:0]  button_pio_external_connection_export,     // button_pio_external_connection.export
		output wire        hps_0_h2f_reset_reset_n,                   //                hps_0_h2f_reset.reset_n
		inout  wire        oc_i2c_master_0_conduit_start_scl_pad_io,  //  oc_i2c_master_0_conduit_start.scl_pad_io
		inout  wire        oc_i2c_master_0_conduit_start_sda_pad_io,  //                               .sda_pad_io
		output wire        clock_bridge_148_5_out_clk_clk,            //     clock_bridge_148_5_out_clk.clk
		output wire        sdram_clk_clk,                             //                      sdram_clk.clk
		output wire [12:0] sdram_wire_addr,                           //                     sdram_wire.addr
		output wire [1:0]  sdram_wire_ba,                             //                               .ba
		output wire        sdram_wire_cas_n,                          //                               .cas_n
		output wire        sdram_wire_cke,                            //                               .cke
		output wire        sdram_wire_cs_n,                           //                               .cs_n
		inout  wire [15:0] sdram_wire_dq,                             //                               .dq
		output wire [1:0]  sdram_wire_dqm,                            //                               .dqm
		output wire        sdram_wire_ras_n,                          //                               .ras_n
		output wire        sdram_wire_we_n,                           //                               .we_n
		input  wire        alt_vip_itc_0_clocked_video_vid_clk,       //    alt_vip_itc_0_clocked_video.vid_clk
		output wire [23:0] alt_vip_itc_0_clocked_video_vid_data,      //                               .vid_data
		output wire        alt_vip_itc_0_clocked_video_underflow,     //                               .underflow
		output wire        alt_vip_itc_0_clocked_video_vid_datavalid, //                               .vid_datavalid
		output wire        alt_vip_itc_0_clocked_video_vid_v_sync,    //                               .vid_v_sync
		output wire        alt_vip_itc_0_clocked_video_vid_h_sync,    //                               .vid_h_sync
		output wire        alt_vip_itc_0_clocked_video_vid_f,         //                               .vid_f
		output wire        alt_vip_itc_0_clocked_video_vid_h,         //                               .vid_h
		output wire        alt_vip_itc_0_clocked_video_vid_v,         //                               .vid_v
		input  wire        clk_clk,                                   //                            clk.clk
		output wire        audio_if_0_conduit_end_XCK,                //         audio_if_0_conduit_end.XCK
		input  wire        audio_if_0_conduit_end_ADCDAT,             //                               .ADCDAT
		input  wire        audio_if_0_conduit_end_ADCLRC,             //                               .ADCLRC
		output wire        audio_if_0_conduit_end_DACDAT,             //                               .DACDAT
		input  wire        audio_if_0_conduit_end_DACLRC,             //                               .DACLRC
		input  wire        audio_if_0_conduit_end_BCLK                //                               .BCLK
	);

	wire          pll_stream_outclk1_clk;                                                                              // pll_stream:outclk_1 -> [LOG_Generate_0:clock, alt_vip_itc_0:is_clk, alt_vip_mix_0:clock, alt_vip_mix_0_control_translator:clk, alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent:clk, alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent_rdata_fifo:clk, alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, alt_vip_tpg_0:clock, alt_vip_vfr_0:clock, alt_vip_vfr_0_avalon_slave_translator:clk, alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent:clk, alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:clk, alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, avalon_st_adapter:in_clk_0_clk, burst_adapter_005:clk, burst_adapter_006:clk, cmd_xbar_mux_007:clk, cmd_xbar_mux_008:clk, crosser:out_clk, crosser_001:out_clk, crosser_003:out_clk, crosser_004:out_clk, crosser_006:in_clk, crosser_007:in_clk, crosser_008:in_clk, crosser_009:in_clk, id_router_007:clk, id_router_008:clk, rsp_xbar_demux_007:clk, rsp_xbar_demux_008:clk, rst_controller_002:clk, timing_adapter_0:clk]
	wire          pll_sdram_outclk1_clk;                                                                               // pll_sdram:outclk_1 -> [addr_router_003:clk, addr_router_004:clk, addr_router_005:clk, alt_vip_vfr_0:master_clock, alt_vip_vfr_0_avalon_master_translator:clk, alt_vip_vfr_0_avalon_master_translator_avalon_universal_master_0_agent:clk, burst_adapter_008:clk, cmd_xbar_demux_003:clk, cmd_xbar_demux_004:clk, cmd_xbar_demux_005:clk, cmd_xbar_mux_010:clk, hps_0:h2f_axi_clk, hps_0_h2f_axi_master_agent:aclk, id_router_010:clk, rsp_xbar_demux_010:clk, rst_controller_001:clk, rst_controller_005:clk, sdram:clk, sdram_s1_translator:clk, sdram_s1_translator_avalon_universal_slave_0_agent:clk, sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:clk, sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, width_adapter_002:clk, width_adapter_003:clk]
	wire          alt_vip_mix_0_dout_endofpacket;                                                                      // alt_vip_mix_0:dout_endofpacket -> alt_vip_itc_0:is_eop
	wire          alt_vip_mix_0_dout_valid;                                                                            // alt_vip_mix_0:dout_valid -> alt_vip_itc_0:is_valid
	wire          alt_vip_mix_0_dout_startofpacket;                                                                    // alt_vip_mix_0:dout_startofpacket -> alt_vip_itc_0:is_sop
	wire   [23:0] alt_vip_mix_0_dout_data;                                                                             // alt_vip_mix_0:dout_data -> alt_vip_itc_0:is_data
	wire          alt_vip_mix_0_dout_ready;                                                                            // alt_vip_itc_0:is_ready -> alt_vip_mix_0:dout_ready
	wire          timing_adapter_0_out_endofpacket;                                                                    // timing_adapter_0:out_endofpacket -> alt_vip_mix_0:din_1_endofpacket
	wire          timing_adapter_0_out_valid;                                                                          // timing_adapter_0:out_valid -> alt_vip_mix_0:din_1_valid
	wire          timing_adapter_0_out_startofpacket;                                                                  // timing_adapter_0:out_startofpacket -> alt_vip_mix_0:din_1_startofpacket
	wire   [23:0] timing_adapter_0_out_data;                                                                           // timing_adapter_0:out_data -> alt_vip_mix_0:din_1_data
	wire          timing_adapter_0_out_ready;                                                                          // alt_vip_mix_0:din_1_ready -> timing_adapter_0:out_ready
	wire          alt_vip_vfr_0_avalon_streaming_source_endofpacket;                                                   // alt_vip_vfr_0:dout_endofpacket -> alt_vip_mix_0:din_2_endofpacket
	wire          alt_vip_vfr_0_avalon_streaming_source_valid;                                                         // alt_vip_vfr_0:dout_valid -> alt_vip_mix_0:din_2_valid
	wire          alt_vip_vfr_0_avalon_streaming_source_startofpacket;                                                 // alt_vip_vfr_0:dout_startofpacket -> alt_vip_mix_0:din_2_startofpacket
	wire   [23:0] alt_vip_vfr_0_avalon_streaming_source_data;                                                          // alt_vip_vfr_0:dout_data -> alt_vip_mix_0:din_2_data
	wire          alt_vip_vfr_0_avalon_streaming_source_ready;                                                         // alt_vip_mix_0:din_2_ready -> alt_vip_vfr_0:dout_ready
	wire          alt_vip_tpg_0_dout_endofpacket;                                                                      // alt_vip_tpg_0:dout_endofpacket -> alt_vip_mix_0:din_0_endofpacket
	wire          alt_vip_tpg_0_dout_valid;                                                                            // alt_vip_tpg_0:dout_valid -> alt_vip_mix_0:din_0_valid
	wire          alt_vip_tpg_0_dout_startofpacket;                                                                    // alt_vip_tpg_0:dout_startofpacket -> alt_vip_mix_0:din_0_startofpacket
	wire   [23:0] alt_vip_tpg_0_dout_data;                                                                             // alt_vip_tpg_0:dout_data -> alt_vip_mix_0:din_0_data
	wire          alt_vip_tpg_0_dout_ready;                                                                            // alt_vip_mix_0:din_0_ready -> alt_vip_tpg_0:dout_ready
	wire          pll_audio_outclk0_clk;                                                                               // pll_audio:outclk_0 -> [AUDIO_IF_0:avs_s1_clk, AUDIO_IF_0_avalon_slave_translator:clk, AUDIO_IF_0_avalon_slave_translator_avalon_universal_slave_0_agent:clk, AUDIO_IF_0_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:clk, AUDIO_IF_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:clk, burst_adapter_007:clk, cmd_xbar_mux_009:clk, crosser_002:out_clk, crosser_005:out_clk, crosser_010:in_clk, crosser_011:in_clk, id_router_009:clk, rsp_xbar_demux_009:clk, rst_controller_003:clk]
	wire          master_secure_master_waitrequest;                                                                    // master_secure_master_translator:av_waitrequest -> master_secure:master_waitrequest
	wire   [31:0] master_secure_master_writedata;                                                                      // master_secure:master_writedata -> master_secure_master_translator:av_writedata
	wire   [31:0] master_secure_master_address;                                                                        // master_secure:master_address -> master_secure_master_translator:av_address
	wire          master_secure_master_write;                                                                          // master_secure:master_write -> master_secure_master_translator:av_write
	wire          master_secure_master_read;                                                                           // master_secure:master_read -> master_secure_master_translator:av_read
	wire   [31:0] master_secure_master_readdata;                                                                       // master_secure_master_translator:av_readdata -> master_secure:master_readdata
	wire    [3:0] master_secure_master_byteenable;                                                                     // master_secure:master_byteenable -> master_secure_master_translator:av_byteenable
	wire          master_secure_master_readdatavalid;                                                                  // master_secure_master_translator:av_readdatavalid -> master_secure:master_readdatavalid
	wire   [31:0] led_pio_s1_translator_avalon_anti_slave_0_writedata;                                                 // led_pio_s1_translator:av_writedata -> led_pio:writedata
	wire    [1:0] led_pio_s1_translator_avalon_anti_slave_0_address;                                                   // led_pio_s1_translator:av_address -> led_pio:address
	wire          led_pio_s1_translator_avalon_anti_slave_0_chipselect;                                                // led_pio_s1_translator:av_chipselect -> led_pio:chipselect
	wire          led_pio_s1_translator_avalon_anti_slave_0_write;                                                     // led_pio_s1_translator:av_write -> led_pio:write_n
	wire   [31:0] led_pio_s1_translator_avalon_anti_slave_0_readdata;                                                  // led_pio:readdata -> led_pio_s1_translator:av_readdata
	wire   [31:0] dipsw_pio_s1_translator_avalon_anti_slave_0_writedata;                                               // dipsw_pio_s1_translator:av_writedata -> dipsw_pio:writedata
	wire    [1:0] dipsw_pio_s1_translator_avalon_anti_slave_0_address;                                                 // dipsw_pio_s1_translator:av_address -> dipsw_pio:address
	wire          dipsw_pio_s1_translator_avalon_anti_slave_0_chipselect;                                              // dipsw_pio_s1_translator:av_chipselect -> dipsw_pio:chipselect
	wire          dipsw_pio_s1_translator_avalon_anti_slave_0_write;                                                   // dipsw_pio_s1_translator:av_write -> dipsw_pio:write_n
	wire   [31:0] dipsw_pio_s1_translator_avalon_anti_slave_0_readdata;                                                // dipsw_pio:readdata -> dipsw_pio_s1_translator:av_readdata
	wire   [31:0] button_pio_s1_translator_avalon_anti_slave_0_writedata;                                              // button_pio_s1_translator:av_writedata -> button_pio:writedata
	wire    [1:0] button_pio_s1_translator_avalon_anti_slave_0_address;                                                // button_pio_s1_translator:av_address -> button_pio:address
	wire          button_pio_s1_translator_avalon_anti_slave_0_chipselect;                                             // button_pio_s1_translator:av_chipselect -> button_pio:chipselect
	wire          button_pio_s1_translator_avalon_anti_slave_0_write;                                                  // button_pio_s1_translator:av_write -> button_pio:write_n
	wire   [31:0] button_pio_s1_translator_avalon_anti_slave_0_readdata;                                               // button_pio:readdata -> button_pio_s1_translator:av_readdata
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest;                              // jtag_uart:av_waitrequest -> jtag_uart_avalon_jtag_slave_translator:av_waitrequest
	wire   [31:0] jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata;                                // jtag_uart_avalon_jtag_slave_translator:av_writedata -> jtag_uart:av_writedata
	wire    [0:0] jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_address;                                  // jtag_uart_avalon_jtag_slave_translator:av_address -> jtag_uart:av_address
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect;                               // jtag_uart_avalon_jtag_slave_translator:av_chipselect -> jtag_uart:av_chipselect
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write;                                    // jtag_uart_avalon_jtag_slave_translator:av_write -> jtag_uart:av_write_n
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read;                                     // jtag_uart_avalon_jtag_slave_translator:av_read -> jtag_uart:av_read_n
	wire   [31:0] jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata;                                 // jtag_uart:av_readdata -> jtag_uart_avalon_jtag_slave_translator:av_readdata
	wire          oc_i2c_master_0_avalon_slave_0_translator_avalon_anti_slave_0_waitrequest;                           // oc_i2c_master_0:wb_ack_o -> oc_i2c_master_0_avalon_slave_0_translator:av_waitrequest
	wire   [31:0] oc_i2c_master_0_avalon_slave_0_translator_avalon_anti_slave_0_writedata;                             // oc_i2c_master_0_avalon_slave_0_translator:av_writedata -> oc_i2c_master_0:wb_dat_i
	wire    [2:0] oc_i2c_master_0_avalon_slave_0_translator_avalon_anti_slave_0_address;                               // oc_i2c_master_0_avalon_slave_0_translator:av_address -> oc_i2c_master_0:wb_adr_i
	wire          oc_i2c_master_0_avalon_slave_0_translator_avalon_anti_slave_0_chipselect;                            // oc_i2c_master_0_avalon_slave_0_translator:av_chipselect -> oc_i2c_master_0:wb_stb_i
	wire          oc_i2c_master_0_avalon_slave_0_translator_avalon_anti_slave_0_write;                                 // oc_i2c_master_0_avalon_slave_0_translator:av_write -> oc_i2c_master_0:wb_we_i
	wire   [31:0] oc_i2c_master_0_avalon_slave_0_translator_avalon_anti_slave_0_readdata;                              // oc_i2c_master_0:wb_dat_o -> oc_i2c_master_0_avalon_slave_0_translator:av_readdata
	wire   [15:0] alt_vip_mix_0_control_translator_avalon_anti_slave_0_writedata;                                      // alt_vip_mix_0_control_translator:av_writedata -> alt_vip_mix_0:control_av_writedata
	wire    [5:0] alt_vip_mix_0_control_translator_avalon_anti_slave_0_address;                                        // alt_vip_mix_0_control_translator:av_address -> alt_vip_mix_0:control_av_address
	wire          alt_vip_mix_0_control_translator_avalon_anti_slave_0_chipselect;                                     // alt_vip_mix_0_control_translator:av_chipselect -> alt_vip_mix_0:control_av_chipselect
	wire          alt_vip_mix_0_control_translator_avalon_anti_slave_0_write;                                          // alt_vip_mix_0_control_translator:av_write -> alt_vip_mix_0:control_av_write
	wire   [15:0] alt_vip_mix_0_control_translator_avalon_anti_slave_0_readdata;                                       // alt_vip_mix_0:control_av_readdata -> alt_vip_mix_0_control_translator:av_readdata
	wire   [31:0] alt_vip_vfr_0_avalon_slave_translator_avalon_anti_slave_0_writedata;                                 // alt_vip_vfr_0_avalon_slave_translator:av_writedata -> alt_vip_vfr_0:slave_writedata
	wire    [4:0] alt_vip_vfr_0_avalon_slave_translator_avalon_anti_slave_0_address;                                   // alt_vip_vfr_0_avalon_slave_translator:av_address -> alt_vip_vfr_0:slave_address
	wire          alt_vip_vfr_0_avalon_slave_translator_avalon_anti_slave_0_write;                                     // alt_vip_vfr_0_avalon_slave_translator:av_write -> alt_vip_vfr_0:slave_write
	wire          alt_vip_vfr_0_avalon_slave_translator_avalon_anti_slave_0_read;                                      // alt_vip_vfr_0_avalon_slave_translator:av_read -> alt_vip_vfr_0:slave_read
	wire   [31:0] alt_vip_vfr_0_avalon_slave_translator_avalon_anti_slave_0_readdata;                                  // alt_vip_vfr_0:slave_readdata -> alt_vip_vfr_0_avalon_slave_translator:av_readdata
	wire   [15:0] audio_if_0_avalon_slave_translator_avalon_anti_slave_0_writedata;                                    // AUDIO_IF_0_avalon_slave_translator:av_writedata -> AUDIO_IF_0:avs_s1_writedata
	wire    [2:0] audio_if_0_avalon_slave_translator_avalon_anti_slave_0_address;                                      // AUDIO_IF_0_avalon_slave_translator:av_address -> AUDIO_IF_0:avs_s1_address
	wire          audio_if_0_avalon_slave_translator_avalon_anti_slave_0_write;                                        // AUDIO_IF_0_avalon_slave_translator:av_write -> AUDIO_IF_0:avs_s1_write
	wire          audio_if_0_avalon_slave_translator_avalon_anti_slave_0_read;                                         // AUDIO_IF_0_avalon_slave_translator:av_read -> AUDIO_IF_0:avs_s1_read
	wire   [15:0] audio_if_0_avalon_slave_translator_avalon_anti_slave_0_readdata;                                     // AUDIO_IF_0:avs_s1_readdata -> AUDIO_IF_0_avalon_slave_translator:av_readdata
	wire          alt_vip_vfr_0_avalon_master_waitrequest;                                                             // alt_vip_vfr_0_avalon_master_translator:av_waitrequest -> alt_vip_vfr_0:master_waitrequest
	wire    [6:0] alt_vip_vfr_0_avalon_master_burstcount;                                                              // alt_vip_vfr_0:master_burstcount -> alt_vip_vfr_0_avalon_master_translator:av_burstcount
	wire   [31:0] alt_vip_vfr_0_avalon_master_address;                                                                 // alt_vip_vfr_0:master_address -> alt_vip_vfr_0_avalon_master_translator:av_address
	wire          alt_vip_vfr_0_avalon_master_read;                                                                    // alt_vip_vfr_0:master_read -> alt_vip_vfr_0_avalon_master_translator:av_read
	wire   [31:0] alt_vip_vfr_0_avalon_master_readdata;                                                                // alt_vip_vfr_0_avalon_master_translator:av_readdata -> alt_vip_vfr_0:master_readdata
	wire          alt_vip_vfr_0_avalon_master_readdatavalid;                                                           // alt_vip_vfr_0_avalon_master_translator:av_readdatavalid -> alt_vip_vfr_0:master_readdatavalid
	wire          sdram_s1_translator_avalon_anti_slave_0_waitrequest;                                                 // sdram:za_waitrequest -> sdram_s1_translator:av_waitrequest
	wire   [15:0] sdram_s1_translator_avalon_anti_slave_0_writedata;                                                   // sdram_s1_translator:av_writedata -> sdram:az_data
	wire   [24:0] sdram_s1_translator_avalon_anti_slave_0_address;                                                     // sdram_s1_translator:av_address -> sdram:az_addr
	wire          sdram_s1_translator_avalon_anti_slave_0_chipselect;                                                  // sdram_s1_translator:av_chipselect -> sdram:az_cs
	wire          sdram_s1_translator_avalon_anti_slave_0_write;                                                       // sdram_s1_translator:av_write -> sdram:az_wr_n
	wire          sdram_s1_translator_avalon_anti_slave_0_read;                                                        // sdram_s1_translator:av_read -> sdram:az_rd_n
	wire   [15:0] sdram_s1_translator_avalon_anti_slave_0_readdata;                                                    // sdram:za_data -> sdram_s1_translator:av_readdata
	wire          sdram_s1_translator_avalon_anti_slave_0_readdatavalid;                                               // sdram:za_valid -> sdram_s1_translator:av_readdatavalid
	wire    [1:0] sdram_s1_translator_avalon_anti_slave_0_byteenable;                                                  // sdram_s1_translator:av_byteenable -> sdram:az_be_n
	wire          master_secure_master_translator_avalon_universal_master_0_waitrequest;                               // master_secure_master_translator_avalon_universal_master_0_agent:av_waitrequest -> master_secure_master_translator:uav_waitrequest
	wire    [2:0] master_secure_master_translator_avalon_universal_master_0_burstcount;                                // master_secure_master_translator:uav_burstcount -> master_secure_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] master_secure_master_translator_avalon_universal_master_0_writedata;                                 // master_secure_master_translator:uav_writedata -> master_secure_master_translator_avalon_universal_master_0_agent:av_writedata
	wire   [31:0] master_secure_master_translator_avalon_universal_master_0_address;                                   // master_secure_master_translator:uav_address -> master_secure_master_translator_avalon_universal_master_0_agent:av_address
	wire          master_secure_master_translator_avalon_universal_master_0_lock;                                      // master_secure_master_translator:uav_lock -> master_secure_master_translator_avalon_universal_master_0_agent:av_lock
	wire          master_secure_master_translator_avalon_universal_master_0_write;                                     // master_secure_master_translator:uav_write -> master_secure_master_translator_avalon_universal_master_0_agent:av_write
	wire          master_secure_master_translator_avalon_universal_master_0_read;                                      // master_secure_master_translator:uav_read -> master_secure_master_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] master_secure_master_translator_avalon_universal_master_0_readdata;                                  // master_secure_master_translator_avalon_universal_master_0_agent:av_readdata -> master_secure_master_translator:uav_readdata
	wire          master_secure_master_translator_avalon_universal_master_0_debugaccess;                               // master_secure_master_translator:uav_debugaccess -> master_secure_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] master_secure_master_translator_avalon_universal_master_0_byteenable;                                // master_secure_master_translator:uav_byteenable -> master_secure_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire          master_secure_master_translator_avalon_universal_master_0_readdatavalid;                             // master_secure_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> master_secure_master_translator:uav_readdatavalid
	wire          hps_0_f2h_axi_slave_agent_altera_axi_master_awvalid;                                                 // hps_0_f2h_axi_slave_agent:awvalid -> hps_0:f2h_AWVALID
	wire    [2:0] hps_0_f2h_axi_slave_agent_altera_axi_master_arsize;                                                  // hps_0_f2h_axi_slave_agent:arsize -> hps_0:f2h_ARSIZE
	wire    [1:0] hps_0_f2h_axi_slave_agent_altera_axi_master_arlock;                                                  // hps_0_f2h_axi_slave_agent:arlock -> hps_0:f2h_ARLOCK
	wire    [3:0] hps_0_f2h_axi_slave_agent_altera_axi_master_awcache;                                                 // hps_0_f2h_axi_slave_agent:awcache -> hps_0:f2h_AWCACHE
	wire          hps_0_f2h_axi_slave_agent_altera_axi_master_arready;                                                 // hps_0:f2h_ARREADY -> hps_0_f2h_axi_slave_agent:arready
	wire    [7:0] hps_0_f2h_axi_slave_agent_altera_axi_master_arid;                                                    // hps_0_f2h_axi_slave_agent:arid -> hps_0:f2h_ARID
	wire          hps_0_f2h_axi_slave_agent_altera_axi_master_rready;                                                  // hps_0_f2h_axi_slave_agent:rready -> hps_0:f2h_RREADY
	wire          hps_0_f2h_axi_slave_agent_altera_axi_master_bready;                                                  // hps_0_f2h_axi_slave_agent:bready -> hps_0:f2h_BREADY
	wire    [2:0] hps_0_f2h_axi_slave_agent_altera_axi_master_awsize;                                                  // hps_0_f2h_axi_slave_agent:awsize -> hps_0:f2h_AWSIZE
	wire    [2:0] hps_0_f2h_axi_slave_agent_altera_axi_master_awprot;                                                  // hps_0_f2h_axi_slave_agent:awprot -> hps_0:f2h_AWPROT
	wire          hps_0_f2h_axi_slave_agent_altera_axi_master_arvalid;                                                 // hps_0_f2h_axi_slave_agent:arvalid -> hps_0:f2h_ARVALID
	wire    [2:0] hps_0_f2h_axi_slave_agent_altera_axi_master_arprot;                                                  // hps_0_f2h_axi_slave_agent:arprot -> hps_0:f2h_ARPROT
	wire    [7:0] hps_0_f2h_axi_slave_agent_altera_axi_master_bid;                                                     // hps_0:f2h_BID -> hps_0_f2h_axi_slave_agent:bid
	wire    [3:0] hps_0_f2h_axi_slave_agent_altera_axi_master_arlen;                                                   // hps_0_f2h_axi_slave_agent:arlen -> hps_0:f2h_ARLEN
	wire          hps_0_f2h_axi_slave_agent_altera_axi_master_awready;                                                 // hps_0:f2h_AWREADY -> hps_0_f2h_axi_slave_agent:awready
	wire    [7:0] hps_0_f2h_axi_slave_agent_altera_axi_master_awid;                                                    // hps_0_f2h_axi_slave_agent:awid -> hps_0:f2h_AWID
	wire          hps_0_f2h_axi_slave_agent_altera_axi_master_bvalid;                                                  // hps_0:f2h_BVALID -> hps_0_f2h_axi_slave_agent:bvalid
	wire    [7:0] hps_0_f2h_axi_slave_agent_altera_axi_master_wid;                                                     // hps_0_f2h_axi_slave_agent:wid -> hps_0:f2h_WID
	wire    [1:0] hps_0_f2h_axi_slave_agent_altera_axi_master_awlock;                                                  // hps_0_f2h_axi_slave_agent:awlock -> hps_0:f2h_AWLOCK
	wire    [1:0] hps_0_f2h_axi_slave_agent_altera_axi_master_awburst;                                                 // hps_0_f2h_axi_slave_agent:awburst -> hps_0:f2h_AWBURST
	wire    [1:0] hps_0_f2h_axi_slave_agent_altera_axi_master_bresp;                                                   // hps_0:f2h_BRESP -> hps_0_f2h_axi_slave_agent:bresp
	wire    [4:0] hps_0_f2h_axi_slave_agent_altera_axi_master_aruser;                                                  // hps_0_f2h_axi_slave_agent:aruser -> hps_0:f2h_ARUSER
	wire    [4:0] hps_0_f2h_axi_slave_agent_altera_axi_master_awuser;                                                  // hps_0_f2h_axi_slave_agent:awuser -> hps_0:f2h_AWUSER
	wire    [7:0] hps_0_f2h_axi_slave_agent_altera_axi_master_wstrb;                                                   // hps_0_f2h_axi_slave_agent:wstrb -> hps_0:f2h_WSTRB
	wire          hps_0_f2h_axi_slave_agent_altera_axi_master_rvalid;                                                  // hps_0:f2h_RVALID -> hps_0_f2h_axi_slave_agent:rvalid
	wire    [1:0] hps_0_f2h_axi_slave_agent_altera_axi_master_arburst;                                                 // hps_0_f2h_axi_slave_agent:arburst -> hps_0:f2h_ARBURST
	wire   [63:0] hps_0_f2h_axi_slave_agent_altera_axi_master_wdata;                                                   // hps_0_f2h_axi_slave_agent:wdata -> hps_0:f2h_WDATA
	wire          hps_0_f2h_axi_slave_agent_altera_axi_master_wready;                                                  // hps_0:f2h_WREADY -> hps_0_f2h_axi_slave_agent:wready
	wire   [63:0] hps_0_f2h_axi_slave_agent_altera_axi_master_rdata;                                                   // hps_0:f2h_RDATA -> hps_0_f2h_axi_slave_agent:rdata
	wire   [31:0] hps_0_f2h_axi_slave_agent_altera_axi_master_araddr;                                                  // hps_0_f2h_axi_slave_agent:araddr -> hps_0:f2h_ARADDR
	wire    [3:0] hps_0_f2h_axi_slave_agent_altera_axi_master_arcache;                                                 // hps_0_f2h_axi_slave_agent:arcache -> hps_0:f2h_ARCACHE
	wire    [3:0] hps_0_f2h_axi_slave_agent_altera_axi_master_awlen;                                                   // hps_0_f2h_axi_slave_agent:awlen -> hps_0:f2h_AWLEN
	wire   [31:0] hps_0_f2h_axi_slave_agent_altera_axi_master_awaddr;                                                  // hps_0_f2h_axi_slave_agent:awaddr -> hps_0:f2h_AWADDR
	wire    [7:0] hps_0_f2h_axi_slave_agent_altera_axi_master_rid;                                                     // hps_0:f2h_RID -> hps_0_f2h_axi_slave_agent:rid
	wire          hps_0_f2h_axi_slave_agent_altera_axi_master_wvalid;                                                  // hps_0_f2h_axi_slave_agent:wvalid -> hps_0:f2h_WVALID
	wire    [1:0] hps_0_f2h_axi_slave_agent_altera_axi_master_rresp;                                                   // hps_0:f2h_RRESP -> hps_0_f2h_axi_slave_agent:rresp
	wire          hps_0_f2h_axi_slave_agent_altera_axi_master_wlast;                                                   // hps_0_f2h_axi_slave_agent:wlast -> hps_0:f2h_WLAST
	wire          hps_0_f2h_axi_slave_agent_altera_axi_master_rlast;                                                   // hps_0:f2h_RLAST -> hps_0_f2h_axi_slave_agent:rlast
	wire          hps_0_h2f_lw_axi_master_awvalid;                                                                     // hps_0:h2f_lw_AWVALID -> hps_0_h2f_lw_axi_master_agent:awvalid
	wire    [2:0] hps_0_h2f_lw_axi_master_arsize;                                                                      // hps_0:h2f_lw_ARSIZE -> hps_0_h2f_lw_axi_master_agent:arsize
	wire    [1:0] hps_0_h2f_lw_axi_master_arlock;                                                                      // hps_0:h2f_lw_ARLOCK -> hps_0_h2f_lw_axi_master_agent:arlock
	wire    [3:0] hps_0_h2f_lw_axi_master_awcache;                                                                     // hps_0:h2f_lw_AWCACHE -> hps_0_h2f_lw_axi_master_agent:awcache
	wire          hps_0_h2f_lw_axi_master_arready;                                                                     // hps_0_h2f_lw_axi_master_agent:arready -> hps_0:h2f_lw_ARREADY
	wire   [11:0] hps_0_h2f_lw_axi_master_arid;                                                                        // hps_0:h2f_lw_ARID -> hps_0_h2f_lw_axi_master_agent:arid
	wire          hps_0_h2f_lw_axi_master_rready;                                                                      // hps_0:h2f_lw_RREADY -> hps_0_h2f_lw_axi_master_agent:rready
	wire          hps_0_h2f_lw_axi_master_bready;                                                                      // hps_0:h2f_lw_BREADY -> hps_0_h2f_lw_axi_master_agent:bready
	wire    [2:0] hps_0_h2f_lw_axi_master_awsize;                                                                      // hps_0:h2f_lw_AWSIZE -> hps_0_h2f_lw_axi_master_agent:awsize
	wire    [2:0] hps_0_h2f_lw_axi_master_awprot;                                                                      // hps_0:h2f_lw_AWPROT -> hps_0_h2f_lw_axi_master_agent:awprot
	wire          hps_0_h2f_lw_axi_master_arvalid;                                                                     // hps_0:h2f_lw_ARVALID -> hps_0_h2f_lw_axi_master_agent:arvalid
	wire    [2:0] hps_0_h2f_lw_axi_master_arprot;                                                                      // hps_0:h2f_lw_ARPROT -> hps_0_h2f_lw_axi_master_agent:arprot
	wire   [11:0] hps_0_h2f_lw_axi_master_bid;                                                                         // hps_0_h2f_lw_axi_master_agent:bid -> hps_0:h2f_lw_BID
	wire    [3:0] hps_0_h2f_lw_axi_master_arlen;                                                                       // hps_0:h2f_lw_ARLEN -> hps_0_h2f_lw_axi_master_agent:arlen
	wire          hps_0_h2f_lw_axi_master_awready;                                                                     // hps_0_h2f_lw_axi_master_agent:awready -> hps_0:h2f_lw_AWREADY
	wire   [11:0] hps_0_h2f_lw_axi_master_awid;                                                                        // hps_0:h2f_lw_AWID -> hps_0_h2f_lw_axi_master_agent:awid
	wire          hps_0_h2f_lw_axi_master_bvalid;                                                                      // hps_0_h2f_lw_axi_master_agent:bvalid -> hps_0:h2f_lw_BVALID
	wire   [11:0] hps_0_h2f_lw_axi_master_wid;                                                                         // hps_0:h2f_lw_WID -> hps_0_h2f_lw_axi_master_agent:wid
	wire    [1:0] hps_0_h2f_lw_axi_master_awlock;                                                                      // hps_0:h2f_lw_AWLOCK -> hps_0_h2f_lw_axi_master_agent:awlock
	wire    [1:0] hps_0_h2f_lw_axi_master_awburst;                                                                     // hps_0:h2f_lw_AWBURST -> hps_0_h2f_lw_axi_master_agent:awburst
	wire    [1:0] hps_0_h2f_lw_axi_master_bresp;                                                                       // hps_0_h2f_lw_axi_master_agent:bresp -> hps_0:h2f_lw_BRESP
	wire    [3:0] hps_0_h2f_lw_axi_master_wstrb;                                                                       // hps_0:h2f_lw_WSTRB -> hps_0_h2f_lw_axi_master_agent:wstrb
	wire          hps_0_h2f_lw_axi_master_rvalid;                                                                      // hps_0_h2f_lw_axi_master_agent:rvalid -> hps_0:h2f_lw_RVALID
	wire   [31:0] hps_0_h2f_lw_axi_master_wdata;                                                                       // hps_0:h2f_lw_WDATA -> hps_0_h2f_lw_axi_master_agent:wdata
	wire          hps_0_h2f_lw_axi_master_wready;                                                                      // hps_0_h2f_lw_axi_master_agent:wready -> hps_0:h2f_lw_WREADY
	wire    [1:0] hps_0_h2f_lw_axi_master_arburst;                                                                     // hps_0:h2f_lw_ARBURST -> hps_0_h2f_lw_axi_master_agent:arburst
	wire   [31:0] hps_0_h2f_lw_axi_master_rdata;                                                                       // hps_0_h2f_lw_axi_master_agent:rdata -> hps_0:h2f_lw_RDATA
	wire   [20:0] hps_0_h2f_lw_axi_master_araddr;                                                                      // hps_0:h2f_lw_ARADDR -> hps_0_h2f_lw_axi_master_agent:araddr
	wire    [3:0] hps_0_h2f_lw_axi_master_arcache;                                                                     // hps_0:h2f_lw_ARCACHE -> hps_0_h2f_lw_axi_master_agent:arcache
	wire    [3:0] hps_0_h2f_lw_axi_master_awlen;                                                                       // hps_0:h2f_lw_AWLEN -> hps_0_h2f_lw_axi_master_agent:awlen
	wire   [20:0] hps_0_h2f_lw_axi_master_awaddr;                                                                      // hps_0:h2f_lw_AWADDR -> hps_0_h2f_lw_axi_master_agent:awaddr
	wire   [11:0] hps_0_h2f_lw_axi_master_rid;                                                                         // hps_0_h2f_lw_axi_master_agent:rid -> hps_0:h2f_lw_RID
	wire          hps_0_h2f_lw_axi_master_wvalid;                                                                      // hps_0:h2f_lw_WVALID -> hps_0_h2f_lw_axi_master_agent:wvalid
	wire    [1:0] hps_0_h2f_lw_axi_master_rresp;                                                                       // hps_0_h2f_lw_axi_master_agent:rresp -> hps_0:h2f_lw_RRESP
	wire          hps_0_h2f_lw_axi_master_wlast;                                                                       // hps_0:h2f_lw_WLAST -> hps_0_h2f_lw_axi_master_agent:wlast
	wire          hps_0_h2f_lw_axi_master_rlast;                                                                       // hps_0_h2f_lw_axi_master_agent:rlast -> hps_0:h2f_lw_RLAST
	wire          led_pio_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                 // led_pio_s1_translator:uav_waitrequest -> led_pio_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] led_pio_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                  // led_pio_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> led_pio_s1_translator:uav_burstcount
	wire   [31:0] led_pio_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                   // led_pio_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> led_pio_s1_translator:uav_writedata
	wire   [20:0] led_pio_s1_translator_avalon_universal_slave_0_agent_m0_address;                                     // led_pio_s1_translator_avalon_universal_slave_0_agent:m0_address -> led_pio_s1_translator:uav_address
	wire          led_pio_s1_translator_avalon_universal_slave_0_agent_m0_write;                                       // led_pio_s1_translator_avalon_universal_slave_0_agent:m0_write -> led_pio_s1_translator:uav_write
	wire          led_pio_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                        // led_pio_s1_translator_avalon_universal_slave_0_agent:m0_lock -> led_pio_s1_translator:uav_lock
	wire          led_pio_s1_translator_avalon_universal_slave_0_agent_m0_read;                                        // led_pio_s1_translator_avalon_universal_slave_0_agent:m0_read -> led_pio_s1_translator:uav_read
	wire   [31:0] led_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                    // led_pio_s1_translator:uav_readdata -> led_pio_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          led_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                               // led_pio_s1_translator:uav_readdatavalid -> led_pio_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          led_pio_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                 // led_pio_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> led_pio_s1_translator:uav_debugaccess
	wire    [3:0] led_pio_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                  // led_pio_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> led_pio_s1_translator:uav_byteenable
	wire          led_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                          // led_pio_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          led_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                // led_pio_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          led_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                        // led_pio_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [113:0] led_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                 // led_pio_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          led_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                // led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> led_pio_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                       // led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> led_pio_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                             // led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> led_pio_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                     // led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> led_pio_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [113:0] led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                              // led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> led_pio_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                             // led_pio_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                           // led_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [33:0] led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                            // led_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                           // led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> led_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                           // led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> led_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                            // led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> led_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                           // led_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          dipsw_pio_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                               // dipsw_pio_s1_translator:uav_waitrequest -> dipsw_pio_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] dipsw_pio_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                // dipsw_pio_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> dipsw_pio_s1_translator:uav_burstcount
	wire   [31:0] dipsw_pio_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                 // dipsw_pio_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> dipsw_pio_s1_translator:uav_writedata
	wire   [20:0] dipsw_pio_s1_translator_avalon_universal_slave_0_agent_m0_address;                                   // dipsw_pio_s1_translator_avalon_universal_slave_0_agent:m0_address -> dipsw_pio_s1_translator:uav_address
	wire          dipsw_pio_s1_translator_avalon_universal_slave_0_agent_m0_write;                                     // dipsw_pio_s1_translator_avalon_universal_slave_0_agent:m0_write -> dipsw_pio_s1_translator:uav_write
	wire          dipsw_pio_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                      // dipsw_pio_s1_translator_avalon_universal_slave_0_agent:m0_lock -> dipsw_pio_s1_translator:uav_lock
	wire          dipsw_pio_s1_translator_avalon_universal_slave_0_agent_m0_read;                                      // dipsw_pio_s1_translator_avalon_universal_slave_0_agent:m0_read -> dipsw_pio_s1_translator:uav_read
	wire   [31:0] dipsw_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                  // dipsw_pio_s1_translator:uav_readdata -> dipsw_pio_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          dipsw_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                             // dipsw_pio_s1_translator:uav_readdatavalid -> dipsw_pio_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          dipsw_pio_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                               // dipsw_pio_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> dipsw_pio_s1_translator:uav_debugaccess
	wire    [3:0] dipsw_pio_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                // dipsw_pio_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> dipsw_pio_s1_translator:uav_byteenable
	wire          dipsw_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                        // dipsw_pio_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> dipsw_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          dipsw_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                              // dipsw_pio_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> dipsw_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          dipsw_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                      // dipsw_pio_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> dipsw_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [113:0] dipsw_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                               // dipsw_pio_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> dipsw_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          dipsw_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                              // dipsw_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> dipsw_pio_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          dipsw_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                     // dipsw_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> dipsw_pio_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          dipsw_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                           // dipsw_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> dipsw_pio_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          dipsw_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                   // dipsw_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> dipsw_pio_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [113:0] dipsw_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                            // dipsw_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> dipsw_pio_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          dipsw_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                           // dipsw_pio_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> dipsw_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          dipsw_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                         // dipsw_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> dipsw_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [33:0] dipsw_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                          // dipsw_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> dipsw_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          dipsw_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                         // dipsw_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> dipsw_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          dipsw_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                         // dipsw_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> dipsw_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] dipsw_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                          // dipsw_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> dipsw_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          dipsw_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                         // dipsw_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> dipsw_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          button_pio_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                              // button_pio_s1_translator:uav_waitrequest -> button_pio_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] button_pio_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                               // button_pio_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> button_pio_s1_translator:uav_burstcount
	wire   [31:0] button_pio_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                // button_pio_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> button_pio_s1_translator:uav_writedata
	wire   [20:0] button_pio_s1_translator_avalon_universal_slave_0_agent_m0_address;                                  // button_pio_s1_translator_avalon_universal_slave_0_agent:m0_address -> button_pio_s1_translator:uav_address
	wire          button_pio_s1_translator_avalon_universal_slave_0_agent_m0_write;                                    // button_pio_s1_translator_avalon_universal_slave_0_agent:m0_write -> button_pio_s1_translator:uav_write
	wire          button_pio_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                     // button_pio_s1_translator_avalon_universal_slave_0_agent:m0_lock -> button_pio_s1_translator:uav_lock
	wire          button_pio_s1_translator_avalon_universal_slave_0_agent_m0_read;                                     // button_pio_s1_translator_avalon_universal_slave_0_agent:m0_read -> button_pio_s1_translator:uav_read
	wire   [31:0] button_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                 // button_pio_s1_translator:uav_readdata -> button_pio_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          button_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                            // button_pio_s1_translator:uav_readdatavalid -> button_pio_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          button_pio_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                              // button_pio_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> button_pio_s1_translator:uav_debugaccess
	wire    [3:0] button_pio_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                               // button_pio_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> button_pio_s1_translator:uav_byteenable
	wire          button_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                       // button_pio_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          button_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                             // button_pio_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          button_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                     // button_pio_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [113:0] button_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                              // button_pio_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          button_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                             // button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> button_pio_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                    // button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> button_pio_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                          // button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> button_pio_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                  // button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> button_pio_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [113:0] button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                           // button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> button_pio_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                          // button_pio_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          button_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                        // button_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> button_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [33:0] button_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                         // button_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> button_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          button_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                        // button_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> button_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          button_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                        // button_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> button_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] button_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                         // button_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> button_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          button_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                        // button_pio_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> button_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                // jtag_uart_avalon_jtag_slave_translator:uav_waitrequest -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                 // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> jtag_uart_avalon_jtag_slave_translator:uav_burstcount
	wire   [31:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                  // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> jtag_uart_avalon_jtag_slave_translator:uav_writedata
	wire   [20:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address;                    // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_address -> jtag_uart_avalon_jtag_slave_translator:uav_address
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write;                      // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_write -> jtag_uart_avalon_jtag_slave_translator:uav_write
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock;                       // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_lock -> jtag_uart_avalon_jtag_slave_translator:uav_lock
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read;                       // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_read -> jtag_uart_avalon_jtag_slave_translator:uav_read
	wire   [31:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                   // jtag_uart_avalon_jtag_slave_translator:uav_readdata -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;              // jtag_uart_avalon_jtag_slave_translator:uav_readdatavalid -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> jtag_uart_avalon_jtag_slave_translator:uav_debugaccess
	wire    [3:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                 // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> jtag_uart_avalon_jtag_slave_translator:uav_byteenable
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;         // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;               // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;       // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [113:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;               // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;      // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;            // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;    // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [113:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;             // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;            // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;          // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [33:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;           // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;          // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;          // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;           // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;          // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest;             // oc_i2c_master_0_avalon_slave_0_translator:uav_waitrequest -> oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount;              // oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_burstcount -> oc_i2c_master_0_avalon_slave_0_translator:uav_burstcount
	wire   [31:0] oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata;               // oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_writedata -> oc_i2c_master_0_avalon_slave_0_translator:uav_writedata
	wire   [20:0] oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address;                 // oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_address -> oc_i2c_master_0_avalon_slave_0_translator:uav_address
	wire          oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write;                   // oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_write -> oc_i2c_master_0_avalon_slave_0_translator:uav_write
	wire          oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock;                    // oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_lock -> oc_i2c_master_0_avalon_slave_0_translator:uav_lock
	wire          oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read;                    // oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_read -> oc_i2c_master_0_avalon_slave_0_translator:uav_read
	wire   [31:0] oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata;                // oc_i2c_master_0_avalon_slave_0_translator:uav_readdata -> oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid;           // oc_i2c_master_0_avalon_slave_0_translator:uav_readdatavalid -> oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess;             // oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_debugaccess -> oc_i2c_master_0_avalon_slave_0_translator:uav_debugaccess
	wire    [3:0] oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable;              // oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:m0_byteenable -> oc_i2c_master_0_avalon_slave_0_translator:uav_byteenable
	wire          oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;      // oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid;            // oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_valid -> oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;    // oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [113:0] oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data;             // oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_data -> oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready;            // oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;   // oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;         // oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket; // oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [113:0] oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;          // oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;         // oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rf_sink_ready -> oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;       // oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [33:0] oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;        // oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;       // oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;       // oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;        // oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;       // oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent_m0_waitrequest;                      // alt_vip_mix_0_control_translator:uav_waitrequest -> alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent_m0_burstcount;                       // alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent:m0_burstcount -> alt_vip_mix_0_control_translator:uav_burstcount
	wire   [31:0] alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent_m0_writedata;                        // alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent:m0_writedata -> alt_vip_mix_0_control_translator:uav_writedata
	wire   [20:0] alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent_m0_address;                          // alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent:m0_address -> alt_vip_mix_0_control_translator:uav_address
	wire          alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent_m0_write;                            // alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent:m0_write -> alt_vip_mix_0_control_translator:uav_write
	wire          alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent_m0_lock;                             // alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent:m0_lock -> alt_vip_mix_0_control_translator:uav_lock
	wire          alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent_m0_read;                             // alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent:m0_read -> alt_vip_mix_0_control_translator:uav_read
	wire   [31:0] alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent_m0_readdata;                         // alt_vip_mix_0_control_translator:uav_readdata -> alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                    // alt_vip_mix_0_control_translator:uav_readdatavalid -> alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent_m0_debugaccess;                      // alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent:m0_debugaccess -> alt_vip_mix_0_control_translator:uav_debugaccess
	wire    [3:0] alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent_m0_byteenable;                       // alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent:m0_byteenable -> alt_vip_mix_0_control_translator:uav_byteenable
	wire          alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;               // alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent_rf_source_valid;                     // alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent:rf_source_valid -> alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;             // alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [113:0] alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent_rf_source_data;                      // alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent:rf_source_data -> alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent_rf_source_ready;                     // alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;            // alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                  // alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;          // alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [113:0] alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                   // alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                  // alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent:rf_sink_ready -> alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                // alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [33:0] alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                 // alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                // alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                // alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                 // alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                // alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                 // alt_vip_vfr_0_avalon_slave_translator:uav_waitrequest -> alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                  // alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> alt_vip_vfr_0_avalon_slave_translator:uav_burstcount
	wire   [31:0] alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                   // alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> alt_vip_vfr_0_avalon_slave_translator:uav_writedata
	wire   [20:0] alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_address;                     // alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent:m0_address -> alt_vip_vfr_0_avalon_slave_translator:uav_address
	wire          alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_write;                       // alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent:m0_write -> alt_vip_vfr_0_avalon_slave_translator:uav_write
	wire          alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_lock;                        // alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent:m0_lock -> alt_vip_vfr_0_avalon_slave_translator:uav_lock
	wire          alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_read;                        // alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent:m0_read -> alt_vip_vfr_0_avalon_slave_translator:uav_read
	wire   [31:0] alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                    // alt_vip_vfr_0_avalon_slave_translator:uav_readdata -> alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;               // alt_vip_vfr_0_avalon_slave_translator:uav_readdatavalid -> alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                 // alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> alt_vip_vfr_0_avalon_slave_translator:uav_debugaccess
	wire    [3:0] alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                  // alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> alt_vip_vfr_0_avalon_slave_translator:uav_byteenable
	wire          alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;          // alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                // alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;        // alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [113:0] alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                 // alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                // alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;       // alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;             // alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;     // alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [113:0] alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;              // alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;             // alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;           // alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [33:0] alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;            // alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;           // alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;           // alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;            // alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;           // alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          audio_if_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest;                    // AUDIO_IF_0_avalon_slave_translator:uav_waitrequest -> AUDIO_IF_0_avalon_slave_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [2:0] audio_if_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_burstcount;                     // AUDIO_IF_0_avalon_slave_translator_avalon_universal_slave_0_agent:m0_burstcount -> AUDIO_IF_0_avalon_slave_translator:uav_burstcount
	wire   [31:0] audio_if_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_writedata;                      // AUDIO_IF_0_avalon_slave_translator_avalon_universal_slave_0_agent:m0_writedata -> AUDIO_IF_0_avalon_slave_translator:uav_writedata
	wire   [20:0] audio_if_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_address;                        // AUDIO_IF_0_avalon_slave_translator_avalon_universal_slave_0_agent:m0_address -> AUDIO_IF_0_avalon_slave_translator:uav_address
	wire          audio_if_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_write;                          // AUDIO_IF_0_avalon_slave_translator_avalon_universal_slave_0_agent:m0_write -> AUDIO_IF_0_avalon_slave_translator:uav_write
	wire          audio_if_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_lock;                           // AUDIO_IF_0_avalon_slave_translator_avalon_universal_slave_0_agent:m0_lock -> AUDIO_IF_0_avalon_slave_translator:uav_lock
	wire          audio_if_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_read;                           // AUDIO_IF_0_avalon_slave_translator_avalon_universal_slave_0_agent:m0_read -> AUDIO_IF_0_avalon_slave_translator:uav_read
	wire   [31:0] audio_if_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_readdata;                       // AUDIO_IF_0_avalon_slave_translator:uav_readdata -> AUDIO_IF_0_avalon_slave_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          audio_if_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                  // AUDIO_IF_0_avalon_slave_translator:uav_readdatavalid -> AUDIO_IF_0_avalon_slave_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          audio_if_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess;                    // AUDIO_IF_0_avalon_slave_translator_avalon_universal_slave_0_agent:m0_debugaccess -> AUDIO_IF_0_avalon_slave_translator:uav_debugaccess
	wire    [3:0] audio_if_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_byteenable;                     // AUDIO_IF_0_avalon_slave_translator_avalon_universal_slave_0_agent:m0_byteenable -> AUDIO_IF_0_avalon_slave_translator:uav_byteenable
	wire          audio_if_0_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;             // AUDIO_IF_0_avalon_slave_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> AUDIO_IF_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          audio_if_0_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_valid;                   // AUDIO_IF_0_avalon_slave_translator_avalon_universal_slave_0_agent:rf_source_valid -> AUDIO_IF_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          audio_if_0_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;           // AUDIO_IF_0_avalon_slave_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> AUDIO_IF_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [113:0] audio_if_0_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_data;                    // AUDIO_IF_0_avalon_slave_translator_avalon_universal_slave_0_agent:rf_source_data -> AUDIO_IF_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          audio_if_0_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_ready;                   // AUDIO_IF_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> AUDIO_IF_0_avalon_slave_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          audio_if_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;          // AUDIO_IF_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> AUDIO_IF_0_avalon_slave_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          audio_if_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                // AUDIO_IF_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> AUDIO_IF_0_avalon_slave_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          audio_if_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;        // AUDIO_IF_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> AUDIO_IF_0_avalon_slave_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [113:0] audio_if_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                 // AUDIO_IF_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> AUDIO_IF_0_avalon_slave_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          audio_if_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                // AUDIO_IF_0_avalon_slave_translator_avalon_universal_slave_0_agent:rf_sink_ready -> AUDIO_IF_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          audio_if_0_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;              // AUDIO_IF_0_avalon_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> AUDIO_IF_0_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [33:0] audio_if_0_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;               // AUDIO_IF_0_avalon_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> AUDIO_IF_0_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          audio_if_0_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;              // AUDIO_IF_0_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> AUDIO_IF_0_avalon_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          audio_if_0_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;              // AUDIO_IF_0_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> AUDIO_IF_0_avalon_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [33:0] audio_if_0_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;               // AUDIO_IF_0_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> AUDIO_IF_0_avalon_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          audio_if_0_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;              // AUDIO_IF_0_avalon_slave_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> AUDIO_IF_0_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          hps_0_h2f_axi_master_awvalid;                                                                        // hps_0:h2f_AWVALID -> hps_0_h2f_axi_master_agent:awvalid
	wire    [2:0] hps_0_h2f_axi_master_arsize;                                                                         // hps_0:h2f_ARSIZE -> hps_0_h2f_axi_master_agent:arsize
	wire    [1:0] hps_0_h2f_axi_master_arlock;                                                                         // hps_0:h2f_ARLOCK -> hps_0_h2f_axi_master_agent:arlock
	wire    [3:0] hps_0_h2f_axi_master_awcache;                                                                        // hps_0:h2f_AWCACHE -> hps_0_h2f_axi_master_agent:awcache
	wire          hps_0_h2f_axi_master_arready;                                                                        // hps_0_h2f_axi_master_agent:arready -> hps_0:h2f_ARREADY
	wire   [11:0] hps_0_h2f_axi_master_arid;                                                                           // hps_0:h2f_ARID -> hps_0_h2f_axi_master_agent:arid
	wire          hps_0_h2f_axi_master_rready;                                                                         // hps_0:h2f_RREADY -> hps_0_h2f_axi_master_agent:rready
	wire          hps_0_h2f_axi_master_bready;                                                                         // hps_0:h2f_BREADY -> hps_0_h2f_axi_master_agent:bready
	wire    [2:0] hps_0_h2f_axi_master_awsize;                                                                         // hps_0:h2f_AWSIZE -> hps_0_h2f_axi_master_agent:awsize
	wire    [2:0] hps_0_h2f_axi_master_awprot;                                                                         // hps_0:h2f_AWPROT -> hps_0_h2f_axi_master_agent:awprot
	wire          hps_0_h2f_axi_master_arvalid;                                                                        // hps_0:h2f_ARVALID -> hps_0_h2f_axi_master_agent:arvalid
	wire    [2:0] hps_0_h2f_axi_master_arprot;                                                                         // hps_0:h2f_ARPROT -> hps_0_h2f_axi_master_agent:arprot
	wire   [11:0] hps_0_h2f_axi_master_bid;                                                                            // hps_0_h2f_axi_master_agent:bid -> hps_0:h2f_BID
	wire    [3:0] hps_0_h2f_axi_master_arlen;                                                                          // hps_0:h2f_ARLEN -> hps_0_h2f_axi_master_agent:arlen
	wire          hps_0_h2f_axi_master_awready;                                                                        // hps_0_h2f_axi_master_agent:awready -> hps_0:h2f_AWREADY
	wire   [11:0] hps_0_h2f_axi_master_awid;                                                                           // hps_0:h2f_AWID -> hps_0_h2f_axi_master_agent:awid
	wire          hps_0_h2f_axi_master_bvalid;                                                                         // hps_0_h2f_axi_master_agent:bvalid -> hps_0:h2f_BVALID
	wire   [11:0] hps_0_h2f_axi_master_wid;                                                                            // hps_0:h2f_WID -> hps_0_h2f_axi_master_agent:wid
	wire    [1:0] hps_0_h2f_axi_master_awlock;                                                                         // hps_0:h2f_AWLOCK -> hps_0_h2f_axi_master_agent:awlock
	wire    [1:0] hps_0_h2f_axi_master_awburst;                                                                        // hps_0:h2f_AWBURST -> hps_0_h2f_axi_master_agent:awburst
	wire    [1:0] hps_0_h2f_axi_master_bresp;                                                                          // hps_0_h2f_axi_master_agent:bresp -> hps_0:h2f_BRESP
	wire   [15:0] hps_0_h2f_axi_master_wstrb;                                                                          // hps_0:h2f_WSTRB -> hps_0_h2f_axi_master_agent:wstrb
	wire          hps_0_h2f_axi_master_rvalid;                                                                         // hps_0_h2f_axi_master_agent:rvalid -> hps_0:h2f_RVALID
	wire  [127:0] hps_0_h2f_axi_master_wdata;                                                                          // hps_0:h2f_WDATA -> hps_0_h2f_axi_master_agent:wdata
	wire          hps_0_h2f_axi_master_wready;                                                                         // hps_0_h2f_axi_master_agent:wready -> hps_0:h2f_WREADY
	wire    [1:0] hps_0_h2f_axi_master_arburst;                                                                        // hps_0:h2f_ARBURST -> hps_0_h2f_axi_master_agent:arburst
	wire  [127:0] hps_0_h2f_axi_master_rdata;                                                                          // hps_0_h2f_axi_master_agent:rdata -> hps_0:h2f_RDATA
	wire   [29:0] hps_0_h2f_axi_master_araddr;                                                                         // hps_0:h2f_ARADDR -> hps_0_h2f_axi_master_agent:araddr
	wire    [3:0] hps_0_h2f_axi_master_arcache;                                                                        // hps_0:h2f_ARCACHE -> hps_0_h2f_axi_master_agent:arcache
	wire    [3:0] hps_0_h2f_axi_master_awlen;                                                                          // hps_0:h2f_AWLEN -> hps_0_h2f_axi_master_agent:awlen
	wire   [29:0] hps_0_h2f_axi_master_awaddr;                                                                         // hps_0:h2f_AWADDR -> hps_0_h2f_axi_master_agent:awaddr
	wire   [11:0] hps_0_h2f_axi_master_rid;                                                                            // hps_0_h2f_axi_master_agent:rid -> hps_0:h2f_RID
	wire          hps_0_h2f_axi_master_wvalid;                                                                         // hps_0:h2f_WVALID -> hps_0_h2f_axi_master_agent:wvalid
	wire    [1:0] hps_0_h2f_axi_master_rresp;                                                                          // hps_0_h2f_axi_master_agent:rresp -> hps_0:h2f_RRESP
	wire          hps_0_h2f_axi_master_wlast;                                                                          // hps_0:h2f_WLAST -> hps_0_h2f_axi_master_agent:wlast
	wire          hps_0_h2f_axi_master_rlast;                                                                          // hps_0_h2f_axi_master_agent:rlast -> hps_0:h2f_RLAST
	wire          alt_vip_vfr_0_avalon_master_translator_avalon_universal_master_0_waitrequest;                        // alt_vip_vfr_0_avalon_master_translator_avalon_universal_master_0_agent:av_waitrequest -> alt_vip_vfr_0_avalon_master_translator:uav_waitrequest
	wire    [8:0] alt_vip_vfr_0_avalon_master_translator_avalon_universal_master_0_burstcount;                         // alt_vip_vfr_0_avalon_master_translator:uav_burstcount -> alt_vip_vfr_0_avalon_master_translator_avalon_universal_master_0_agent:av_burstcount
	wire   [31:0] alt_vip_vfr_0_avalon_master_translator_avalon_universal_master_0_writedata;                          // alt_vip_vfr_0_avalon_master_translator:uav_writedata -> alt_vip_vfr_0_avalon_master_translator_avalon_universal_master_0_agent:av_writedata
	wire   [31:0] alt_vip_vfr_0_avalon_master_translator_avalon_universal_master_0_address;                            // alt_vip_vfr_0_avalon_master_translator:uav_address -> alt_vip_vfr_0_avalon_master_translator_avalon_universal_master_0_agent:av_address
	wire          alt_vip_vfr_0_avalon_master_translator_avalon_universal_master_0_lock;                               // alt_vip_vfr_0_avalon_master_translator:uav_lock -> alt_vip_vfr_0_avalon_master_translator_avalon_universal_master_0_agent:av_lock
	wire          alt_vip_vfr_0_avalon_master_translator_avalon_universal_master_0_write;                              // alt_vip_vfr_0_avalon_master_translator:uav_write -> alt_vip_vfr_0_avalon_master_translator_avalon_universal_master_0_agent:av_write
	wire          alt_vip_vfr_0_avalon_master_translator_avalon_universal_master_0_read;                               // alt_vip_vfr_0_avalon_master_translator:uav_read -> alt_vip_vfr_0_avalon_master_translator_avalon_universal_master_0_agent:av_read
	wire   [31:0] alt_vip_vfr_0_avalon_master_translator_avalon_universal_master_0_readdata;                           // alt_vip_vfr_0_avalon_master_translator_avalon_universal_master_0_agent:av_readdata -> alt_vip_vfr_0_avalon_master_translator:uav_readdata
	wire          alt_vip_vfr_0_avalon_master_translator_avalon_universal_master_0_debugaccess;                        // alt_vip_vfr_0_avalon_master_translator:uav_debugaccess -> alt_vip_vfr_0_avalon_master_translator_avalon_universal_master_0_agent:av_debugaccess
	wire    [3:0] alt_vip_vfr_0_avalon_master_translator_avalon_universal_master_0_byteenable;                         // alt_vip_vfr_0_avalon_master_translator:uav_byteenable -> alt_vip_vfr_0_avalon_master_translator_avalon_universal_master_0_agent:av_byteenable
	wire          alt_vip_vfr_0_avalon_master_translator_avalon_universal_master_0_readdatavalid;                      // alt_vip_vfr_0_avalon_master_translator_avalon_universal_master_0_agent:av_readdatavalid -> alt_vip_vfr_0_avalon_master_translator:uav_readdatavalid
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest;                                   // sdram_s1_translator:uav_waitrequest -> sdram_s1_translator_avalon_universal_slave_0_agent:m0_waitrequest
	wire    [1:0] sdram_s1_translator_avalon_universal_slave_0_agent_m0_burstcount;                                    // sdram_s1_translator_avalon_universal_slave_0_agent:m0_burstcount -> sdram_s1_translator:uav_burstcount
	wire   [15:0] sdram_s1_translator_avalon_universal_slave_0_agent_m0_writedata;                                     // sdram_s1_translator_avalon_universal_slave_0_agent:m0_writedata -> sdram_s1_translator:uav_writedata
	wire   [31:0] sdram_s1_translator_avalon_universal_slave_0_agent_m0_address;                                       // sdram_s1_translator_avalon_universal_slave_0_agent:m0_address -> sdram_s1_translator:uav_address
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_m0_write;                                         // sdram_s1_translator_avalon_universal_slave_0_agent:m0_write -> sdram_s1_translator:uav_write
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_m0_lock;                                          // sdram_s1_translator_avalon_universal_slave_0_agent:m0_lock -> sdram_s1_translator:uav_lock
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_m0_read;                                          // sdram_s1_translator_avalon_universal_slave_0_agent:m0_read -> sdram_s1_translator:uav_read
	wire   [15:0] sdram_s1_translator_avalon_universal_slave_0_agent_m0_readdata;                                      // sdram_s1_translator:uav_readdata -> sdram_s1_translator_avalon_universal_slave_0_agent:m0_readdata
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid;                                 // sdram_s1_translator:uav_readdatavalid -> sdram_s1_translator_avalon_universal_slave_0_agent:m0_readdatavalid
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess;                                   // sdram_s1_translator_avalon_universal_slave_0_agent:m0_debugaccess -> sdram_s1_translator:uav_debugaccess
	wire    [1:0] sdram_s1_translator_avalon_universal_slave_0_agent_m0_byteenable;                                    // sdram_s1_translator_avalon_universal_slave_0_agent:m0_byteenable -> sdram_s1_translator:uav_byteenable
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket;                            // sdram_s1_translator_avalon_universal_slave_0_agent:rf_source_endofpacket -> sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_endofpacket
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_valid;                                  // sdram_s1_translator_avalon_universal_slave_0_agent:rf_source_valid -> sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_valid
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket;                          // sdram_s1_translator_avalon_universal_slave_0_agent:rf_source_startofpacket -> sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_startofpacket
	wire  [108:0] sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_data;                                   // sdram_s1_translator_avalon_universal_slave_0_agent:rf_source_data -> sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_data
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_ready;                                  // sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:in_ready -> sdram_s1_translator_avalon_universal_slave_0_agent:rf_source_ready
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket;                         // sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_endofpacket -> sdram_s1_translator_avalon_universal_slave_0_agent:rf_sink_endofpacket
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid;                               // sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_valid -> sdram_s1_translator_avalon_universal_slave_0_agent:rf_sink_valid
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket;                       // sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_startofpacket -> sdram_s1_translator_avalon_universal_slave_0_agent:rf_sink_startofpacket
	wire  [108:0] sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data;                                // sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_data -> sdram_s1_translator_avalon_universal_slave_0_agent:rf_sink_data
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready;                               // sdram_s1_translator_avalon_universal_slave_0_agent:rf_sink_ready -> sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:out_ready
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid;                             // sdram_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_valid -> sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_valid
	wire   [17:0] sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data;                              // sdram_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_data -> sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_data
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready;                             // sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:in_ready -> sdram_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_src_ready
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid;                             // sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_valid -> sdram_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_valid
	wire   [17:0] sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data;                              // sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_data -> sdram_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_data
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready;                             // sdram_s1_translator_avalon_universal_slave_0_agent:rdata_fifo_sink_ready -> sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:out_ready
	wire          master_secure_master_translator_avalon_universal_master_0_agent_cp_endofpacket;                      // master_secure_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router:sink_endofpacket
	wire          master_secure_master_translator_avalon_universal_master_0_agent_cp_valid;                            // master_secure_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router:sink_valid
	wire          master_secure_master_translator_avalon_universal_master_0_agent_cp_startofpacket;                    // master_secure_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router:sink_startofpacket
	wire  [114:0] master_secure_master_translator_avalon_universal_master_0_agent_cp_data;                             // master_secure_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router:sink_data
	wire          master_secure_master_translator_avalon_universal_master_0_agent_cp_ready;                            // addr_router:sink_ready -> master_secure_master_translator_avalon_universal_master_0_agent:cp_ready
	wire          hps_0_f2h_axi_slave_agent_write_rp_endofpacket;                                                      // hps_0_f2h_axi_slave_agent:write_rp_endofpacket -> id_router:sink_endofpacket
	wire          hps_0_f2h_axi_slave_agent_write_rp_valid;                                                            // hps_0_f2h_axi_slave_agent:write_rp_valid -> id_router:sink_valid
	wire          hps_0_f2h_axi_slave_agent_write_rp_startofpacket;                                                    // hps_0_f2h_axi_slave_agent:write_rp_startofpacket -> id_router:sink_startofpacket
	wire  [150:0] hps_0_f2h_axi_slave_agent_write_rp_data;                                                             // hps_0_f2h_axi_slave_agent:write_rp_data -> id_router:sink_data
	wire          hps_0_f2h_axi_slave_agent_write_rp_ready;                                                            // id_router:sink_ready -> hps_0_f2h_axi_slave_agent:write_rp_ready
	wire          hps_0_f2h_axi_slave_agent_read_rp_endofpacket;                                                       // hps_0_f2h_axi_slave_agent:read_rp_endofpacket -> id_router_001:sink_endofpacket
	wire          hps_0_f2h_axi_slave_agent_read_rp_valid;                                                             // hps_0_f2h_axi_slave_agent:read_rp_valid -> id_router_001:sink_valid
	wire          hps_0_f2h_axi_slave_agent_read_rp_startofpacket;                                                     // hps_0_f2h_axi_slave_agent:read_rp_startofpacket -> id_router_001:sink_startofpacket
	wire  [150:0] hps_0_f2h_axi_slave_agent_read_rp_data;                                                              // hps_0_f2h_axi_slave_agent:read_rp_data -> id_router_001:sink_data
	wire          hps_0_f2h_axi_slave_agent_read_rp_ready;                                                             // id_router_001:sink_ready -> hps_0_f2h_axi_slave_agent:read_rp_ready
	wire          hps_0_h2f_lw_axi_master_agent_write_cp_endofpacket;                                                  // hps_0_h2f_lw_axi_master_agent:write_cp_endofpacket -> addr_router_001:sink_endofpacket
	wire          hps_0_h2f_lw_axi_master_agent_write_cp_valid;                                                        // hps_0_h2f_lw_axi_master_agent:write_cp_valid -> addr_router_001:sink_valid
	wire          hps_0_h2f_lw_axi_master_agent_write_cp_startofpacket;                                                // hps_0_h2f_lw_axi_master_agent:write_cp_startofpacket -> addr_router_001:sink_startofpacket
	wire  [112:0] hps_0_h2f_lw_axi_master_agent_write_cp_data;                                                         // hps_0_h2f_lw_axi_master_agent:write_cp_data -> addr_router_001:sink_data
	wire          hps_0_h2f_lw_axi_master_agent_write_cp_ready;                                                        // addr_router_001:sink_ready -> hps_0_h2f_lw_axi_master_agent:write_cp_ready
	wire          hps_0_h2f_lw_axi_master_agent_read_cp_endofpacket;                                                   // hps_0_h2f_lw_axi_master_agent:read_cp_endofpacket -> addr_router_002:sink_endofpacket
	wire          hps_0_h2f_lw_axi_master_agent_read_cp_valid;                                                         // hps_0_h2f_lw_axi_master_agent:read_cp_valid -> addr_router_002:sink_valid
	wire          hps_0_h2f_lw_axi_master_agent_read_cp_startofpacket;                                                 // hps_0_h2f_lw_axi_master_agent:read_cp_startofpacket -> addr_router_002:sink_startofpacket
	wire  [112:0] hps_0_h2f_lw_axi_master_agent_read_cp_data;                                                          // hps_0_h2f_lw_axi_master_agent:read_cp_data -> addr_router_002:sink_data
	wire          hps_0_h2f_lw_axi_master_agent_read_cp_ready;                                                         // addr_router_002:sink_ready -> hps_0_h2f_lw_axi_master_agent:read_cp_ready
	wire          led_pio_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                 // led_pio_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_002:sink_endofpacket
	wire          led_pio_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                       // led_pio_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_002:sink_valid
	wire          led_pio_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                               // led_pio_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_002:sink_startofpacket
	wire  [112:0] led_pio_s1_translator_avalon_universal_slave_0_agent_rp_data;                                        // led_pio_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_002:sink_data
	wire          led_pio_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                       // id_router_002:sink_ready -> led_pio_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          dipsw_pio_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                               // dipsw_pio_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_003:sink_endofpacket
	wire          dipsw_pio_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                     // dipsw_pio_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_003:sink_valid
	wire          dipsw_pio_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                             // dipsw_pio_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_003:sink_startofpacket
	wire  [112:0] dipsw_pio_s1_translator_avalon_universal_slave_0_agent_rp_data;                                      // dipsw_pio_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_003:sink_data
	wire          dipsw_pio_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                     // id_router_003:sink_ready -> dipsw_pio_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          button_pio_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                              // button_pio_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_004:sink_endofpacket
	wire          button_pio_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                    // button_pio_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_004:sink_valid
	wire          button_pio_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                            // button_pio_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_004:sink_startofpacket
	wire  [112:0] button_pio_s1_translator_avalon_universal_slave_0_agent_rp_data;                                     // button_pio_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_004:sink_data
	wire          button_pio_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                    // id_router_004:sink_ready -> button_pio_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_005:sink_endofpacket
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid;                      // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_005:sink_valid
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;              // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_005:sink_startofpacket
	wire  [112:0] jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data;                       // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_005:sink_data
	wire          jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready;                      // id_router_005:sink_ready -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket;             // oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_006:sink_endofpacket
	wire          oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid;                   // oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_006:sink_valid
	wire          oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket;           // oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_006:sink_startofpacket
	wire  [112:0] oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data;                    // oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_data -> id_router_006:sink_data
	wire          oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready;                   // id_router_006:sink_ready -> oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:rp_ready
	wire          alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent_rp_endofpacket;                      // alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_007:sink_endofpacket
	wire          alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent_rp_valid;                            // alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_007:sink_valid
	wire          alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent_rp_startofpacket;                    // alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_007:sink_startofpacket
	wire  [112:0] alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent_rp_data;                             // alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent:rp_data -> id_router_007:sink_data
	wire          alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent_rp_ready;                            // id_router_007:sink_ready -> alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent:rp_ready
	wire          alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                 // alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_008:sink_endofpacket
	wire          alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent_rp_valid;                       // alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_008:sink_valid
	wire          alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;               // alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_008:sink_startofpacket
	wire  [112:0] alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent_rp_data;                        // alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_008:sink_data
	wire          alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent_rp_ready;                       // id_router_008:sink_ready -> alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          audio_if_0_avalon_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket;                    // AUDIO_IF_0_avalon_slave_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_009:sink_endofpacket
	wire          audio_if_0_avalon_slave_translator_avalon_universal_slave_0_agent_rp_valid;                          // AUDIO_IF_0_avalon_slave_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_009:sink_valid
	wire          audio_if_0_avalon_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket;                  // AUDIO_IF_0_avalon_slave_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_009:sink_startofpacket
	wire  [112:0] audio_if_0_avalon_slave_translator_avalon_universal_slave_0_agent_rp_data;                           // AUDIO_IF_0_avalon_slave_translator_avalon_universal_slave_0_agent:rp_data -> id_router_009:sink_data
	wire          audio_if_0_avalon_slave_translator_avalon_universal_slave_0_agent_rp_ready;                          // id_router_009:sink_ready -> AUDIO_IF_0_avalon_slave_translator_avalon_universal_slave_0_agent:rp_ready
	wire          hps_0_h2f_axi_master_agent_write_cp_endofpacket;                                                     // hps_0_h2f_axi_master_agent:write_cp_endofpacket -> addr_router_003:sink_endofpacket
	wire          hps_0_h2f_axi_master_agent_write_cp_valid;                                                           // hps_0_h2f_axi_master_agent:write_cp_valid -> addr_router_003:sink_valid
	wire          hps_0_h2f_axi_master_agent_write_cp_startofpacket;                                                   // hps_0_h2f_axi_master_agent:write_cp_startofpacket -> addr_router_003:sink_startofpacket
	wire  [233:0] hps_0_h2f_axi_master_agent_write_cp_data;                                                            // hps_0_h2f_axi_master_agent:write_cp_data -> addr_router_003:sink_data
	wire          hps_0_h2f_axi_master_agent_write_cp_ready;                                                           // addr_router_003:sink_ready -> hps_0_h2f_axi_master_agent:write_cp_ready
	wire          hps_0_h2f_axi_master_agent_read_cp_endofpacket;                                                      // hps_0_h2f_axi_master_agent:read_cp_endofpacket -> addr_router_004:sink_endofpacket
	wire          hps_0_h2f_axi_master_agent_read_cp_valid;                                                            // hps_0_h2f_axi_master_agent:read_cp_valid -> addr_router_004:sink_valid
	wire          hps_0_h2f_axi_master_agent_read_cp_startofpacket;                                                    // hps_0_h2f_axi_master_agent:read_cp_startofpacket -> addr_router_004:sink_startofpacket
	wire  [233:0] hps_0_h2f_axi_master_agent_read_cp_data;                                                             // hps_0_h2f_axi_master_agent:read_cp_data -> addr_router_004:sink_data
	wire          hps_0_h2f_axi_master_agent_read_cp_ready;                                                            // addr_router_004:sink_ready -> hps_0_h2f_axi_master_agent:read_cp_ready
	wire          alt_vip_vfr_0_avalon_master_translator_avalon_universal_master_0_agent_cp_endofpacket;               // alt_vip_vfr_0_avalon_master_translator_avalon_universal_master_0_agent:cp_endofpacket -> addr_router_005:sink_endofpacket
	wire          alt_vip_vfr_0_avalon_master_translator_avalon_universal_master_0_agent_cp_valid;                     // alt_vip_vfr_0_avalon_master_translator_avalon_universal_master_0_agent:cp_valid -> addr_router_005:sink_valid
	wire          alt_vip_vfr_0_avalon_master_translator_avalon_universal_master_0_agent_cp_startofpacket;             // alt_vip_vfr_0_avalon_master_translator_avalon_universal_master_0_agent:cp_startofpacket -> addr_router_005:sink_startofpacket
	wire  [125:0] alt_vip_vfr_0_avalon_master_translator_avalon_universal_master_0_agent_cp_data;                      // alt_vip_vfr_0_avalon_master_translator_avalon_universal_master_0_agent:cp_data -> addr_router_005:sink_data
	wire          alt_vip_vfr_0_avalon_master_translator_avalon_universal_master_0_agent_cp_ready;                     // addr_router_005:sink_ready -> alt_vip_vfr_0_avalon_master_translator_avalon_universal_master_0_agent:cp_ready
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket;                                   // sdram_s1_translator_avalon_universal_slave_0_agent:rp_endofpacket -> id_router_010:sink_endofpacket
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rp_valid;                                         // sdram_s1_translator_avalon_universal_slave_0_agent:rp_valid -> id_router_010:sink_valid
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket;                                 // sdram_s1_translator_avalon_universal_slave_0_agent:rp_startofpacket -> id_router_010:sink_startofpacket
	wire  [107:0] sdram_s1_translator_avalon_universal_slave_0_agent_rp_data;                                          // sdram_s1_translator_avalon_universal_slave_0_agent:rp_data -> id_router_010:sink_data
	wire          sdram_s1_translator_avalon_universal_slave_0_agent_rp_ready;                                         // id_router_010:sink_ready -> sdram_s1_translator_avalon_universal_slave_0_agent:rp_ready
	wire          addr_router_src_endofpacket;                                                                         // addr_router:src_endofpacket -> limiter:cmd_sink_endofpacket
	wire          addr_router_src_valid;                                                                               // addr_router:src_valid -> limiter:cmd_sink_valid
	wire          addr_router_src_startofpacket;                                                                       // addr_router:src_startofpacket -> limiter:cmd_sink_startofpacket
	wire  [114:0] addr_router_src_data;                                                                                // addr_router:src_data -> limiter:cmd_sink_data
	wire    [1:0] addr_router_src_channel;                                                                             // addr_router:src_channel -> limiter:cmd_sink_channel
	wire          addr_router_src_ready;                                                                               // limiter:cmd_sink_ready -> addr_router:src_ready
	wire          limiter_rsp_src_endofpacket;                                                                         // limiter:rsp_src_endofpacket -> master_secure_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          limiter_rsp_src_valid;                                                                               // limiter:rsp_src_valid -> master_secure_master_translator_avalon_universal_master_0_agent:rp_valid
	wire          limiter_rsp_src_startofpacket;                                                                       // limiter:rsp_src_startofpacket -> master_secure_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [114:0] limiter_rsp_src_data;                                                                                // limiter:rsp_src_data -> master_secure_master_translator_avalon_universal_master_0_agent:rp_data
	wire    [1:0] limiter_rsp_src_channel;                                                                             // limiter:rsp_src_channel -> master_secure_master_translator_avalon_universal_master_0_agent:rp_channel
	wire          limiter_rsp_src_ready;                                                                               // master_secure_master_translator_avalon_universal_master_0_agent:rp_ready -> limiter:rsp_src_ready
	wire          addr_router_001_src_endofpacket;                                                                     // addr_router_001:src_endofpacket -> limiter_001:cmd_sink_endofpacket
	wire          addr_router_001_src_valid;                                                                           // addr_router_001:src_valid -> limiter_001:cmd_sink_valid
	wire          addr_router_001_src_startofpacket;                                                                   // addr_router_001:src_startofpacket -> limiter_001:cmd_sink_startofpacket
	wire  [112:0] addr_router_001_src_data;                                                                            // addr_router_001:src_data -> limiter_001:cmd_sink_data
	wire    [7:0] addr_router_001_src_channel;                                                                         // addr_router_001:src_channel -> limiter_001:cmd_sink_channel
	wire          addr_router_001_src_ready;                                                                           // limiter_001:cmd_sink_ready -> addr_router_001:src_ready
	wire          limiter_001_rsp_src_endofpacket;                                                                     // limiter_001:rsp_src_endofpacket -> hps_0_h2f_lw_axi_master_agent:write_rp_endofpacket
	wire          limiter_001_rsp_src_valid;                                                                           // limiter_001:rsp_src_valid -> hps_0_h2f_lw_axi_master_agent:write_rp_valid
	wire          limiter_001_rsp_src_startofpacket;                                                                   // limiter_001:rsp_src_startofpacket -> hps_0_h2f_lw_axi_master_agent:write_rp_startofpacket
	wire  [112:0] limiter_001_rsp_src_data;                                                                            // limiter_001:rsp_src_data -> hps_0_h2f_lw_axi_master_agent:write_rp_data
	wire    [7:0] limiter_001_rsp_src_channel;                                                                         // limiter_001:rsp_src_channel -> hps_0_h2f_lw_axi_master_agent:write_rp_channel
	wire          limiter_001_rsp_src_ready;                                                                           // hps_0_h2f_lw_axi_master_agent:write_rp_ready -> limiter_001:rsp_src_ready
	wire          addr_router_002_src_endofpacket;                                                                     // addr_router_002:src_endofpacket -> limiter_002:cmd_sink_endofpacket
	wire          addr_router_002_src_valid;                                                                           // addr_router_002:src_valid -> limiter_002:cmd_sink_valid
	wire          addr_router_002_src_startofpacket;                                                                   // addr_router_002:src_startofpacket -> limiter_002:cmd_sink_startofpacket
	wire  [112:0] addr_router_002_src_data;                                                                            // addr_router_002:src_data -> limiter_002:cmd_sink_data
	wire    [7:0] addr_router_002_src_channel;                                                                         // addr_router_002:src_channel -> limiter_002:cmd_sink_channel
	wire          addr_router_002_src_ready;                                                                           // limiter_002:cmd_sink_ready -> addr_router_002:src_ready
	wire          limiter_002_rsp_src_endofpacket;                                                                     // limiter_002:rsp_src_endofpacket -> hps_0_h2f_lw_axi_master_agent:read_rp_endofpacket
	wire          limiter_002_rsp_src_valid;                                                                           // limiter_002:rsp_src_valid -> hps_0_h2f_lw_axi_master_agent:read_rp_valid
	wire          limiter_002_rsp_src_startofpacket;                                                                   // limiter_002:rsp_src_startofpacket -> hps_0_h2f_lw_axi_master_agent:read_rp_startofpacket
	wire  [112:0] limiter_002_rsp_src_data;                                                                            // limiter_002:rsp_src_data -> hps_0_h2f_lw_axi_master_agent:read_rp_data
	wire    [7:0] limiter_002_rsp_src_channel;                                                                         // limiter_002:rsp_src_channel -> hps_0_h2f_lw_axi_master_agent:read_rp_channel
	wire          limiter_002_rsp_src_ready;                                                                           // hps_0_h2f_lw_axi_master_agent:read_rp_ready -> limiter_002:rsp_src_ready
	wire          burst_adapter_source0_endofpacket;                                                                   // burst_adapter:source0_endofpacket -> led_pio_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          burst_adapter_source0_valid;                                                                         // burst_adapter:source0_valid -> led_pio_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          burst_adapter_source0_startofpacket;                                                                 // burst_adapter:source0_startofpacket -> led_pio_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [112:0] burst_adapter_source0_data;                                                                          // burst_adapter:source0_data -> led_pio_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire          burst_adapter_source0_ready;                                                                         // led_pio_s1_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter:source0_ready
	wire    [7:0] burst_adapter_source0_channel;                                                                       // burst_adapter:source0_channel -> led_pio_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          burst_adapter_001_source0_endofpacket;                                                               // burst_adapter_001:source0_endofpacket -> dipsw_pio_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          burst_adapter_001_source0_valid;                                                                     // burst_adapter_001:source0_valid -> dipsw_pio_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          burst_adapter_001_source0_startofpacket;                                                             // burst_adapter_001:source0_startofpacket -> dipsw_pio_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [112:0] burst_adapter_001_source0_data;                                                                      // burst_adapter_001:source0_data -> dipsw_pio_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire          burst_adapter_001_source0_ready;                                                                     // dipsw_pio_s1_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_001:source0_ready
	wire    [7:0] burst_adapter_001_source0_channel;                                                                   // burst_adapter_001:source0_channel -> dipsw_pio_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          burst_adapter_002_source0_endofpacket;                                                               // burst_adapter_002:source0_endofpacket -> button_pio_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          burst_adapter_002_source0_valid;                                                                     // burst_adapter_002:source0_valid -> button_pio_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          burst_adapter_002_source0_startofpacket;                                                             // burst_adapter_002:source0_startofpacket -> button_pio_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [112:0] burst_adapter_002_source0_data;                                                                      // burst_adapter_002:source0_data -> button_pio_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire          burst_adapter_002_source0_ready;                                                                     // button_pio_s1_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_002:source0_ready
	wire    [7:0] burst_adapter_002_source0_channel;                                                                   // burst_adapter_002:source0_channel -> button_pio_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          burst_adapter_003_source0_endofpacket;                                                               // burst_adapter_003:source0_endofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          burst_adapter_003_source0_valid;                                                                     // burst_adapter_003:source0_valid -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          burst_adapter_003_source0_startofpacket;                                                             // burst_adapter_003:source0_startofpacket -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [112:0] burst_adapter_003_source0_data;                                                                      // burst_adapter_003:source0_data -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire          burst_adapter_003_source0_ready;                                                                     // jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_003:source0_ready
	wire    [7:0] burst_adapter_003_source0_channel;                                                                   // burst_adapter_003:source0_channel -> jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          burst_adapter_004_source0_endofpacket;                                                               // burst_adapter_004:source0_endofpacket -> oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          burst_adapter_004_source0_valid;                                                                     // burst_adapter_004:source0_valid -> oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_valid
	wire          burst_adapter_004_source0_startofpacket;                                                             // burst_adapter_004:source0_startofpacket -> oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [112:0] burst_adapter_004_source0_data;                                                                      // burst_adapter_004:source0_data -> oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_data
	wire          burst_adapter_004_source0_ready;                                                                     // oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_004:source0_ready
	wire    [7:0] burst_adapter_004_source0_channel;                                                                   // burst_adapter_004:source0_channel -> oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:cp_channel
	wire          burst_adapter_005_source0_endofpacket;                                                               // burst_adapter_005:source0_endofpacket -> alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          burst_adapter_005_source0_valid;                                                                     // burst_adapter_005:source0_valid -> alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent:cp_valid
	wire          burst_adapter_005_source0_startofpacket;                                                             // burst_adapter_005:source0_startofpacket -> alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [112:0] burst_adapter_005_source0_data;                                                                      // burst_adapter_005:source0_data -> alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent:cp_data
	wire          burst_adapter_005_source0_ready;                                                                     // alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_005:source0_ready
	wire    [7:0] burst_adapter_005_source0_channel;                                                                   // burst_adapter_005:source0_channel -> alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent:cp_channel
	wire          burst_adapter_006_source0_endofpacket;                                                               // burst_adapter_006:source0_endofpacket -> alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          burst_adapter_006_source0_valid;                                                                     // burst_adapter_006:source0_valid -> alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          burst_adapter_006_source0_startofpacket;                                                             // burst_adapter_006:source0_startofpacket -> alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [112:0] burst_adapter_006_source0_data;                                                                      // burst_adapter_006:source0_data -> alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire          burst_adapter_006_source0_ready;                                                                     // alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_006:source0_ready
	wire    [7:0] burst_adapter_006_source0_channel;                                                                   // burst_adapter_006:source0_channel -> alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          burst_adapter_007_source0_endofpacket;                                                               // burst_adapter_007:source0_endofpacket -> AUDIO_IF_0_avalon_slave_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          burst_adapter_007_source0_valid;                                                                     // burst_adapter_007:source0_valid -> AUDIO_IF_0_avalon_slave_translator_avalon_universal_slave_0_agent:cp_valid
	wire          burst_adapter_007_source0_startofpacket;                                                             // burst_adapter_007:source0_startofpacket -> AUDIO_IF_0_avalon_slave_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [112:0] burst_adapter_007_source0_data;                                                                      // burst_adapter_007:source0_data -> AUDIO_IF_0_avalon_slave_translator_avalon_universal_slave_0_agent:cp_data
	wire          burst_adapter_007_source0_ready;                                                                     // AUDIO_IF_0_avalon_slave_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_007:source0_ready
	wire    [7:0] burst_adapter_007_source0_channel;                                                                   // burst_adapter_007:source0_channel -> AUDIO_IF_0_avalon_slave_translator_avalon_universal_slave_0_agent:cp_channel
	wire          burst_adapter_008_source0_endofpacket;                                                               // burst_adapter_008:source0_endofpacket -> sdram_s1_translator_avalon_universal_slave_0_agent:cp_endofpacket
	wire          burst_adapter_008_source0_valid;                                                                     // burst_adapter_008:source0_valid -> sdram_s1_translator_avalon_universal_slave_0_agent:cp_valid
	wire          burst_adapter_008_source0_startofpacket;                                                             // burst_adapter_008:source0_startofpacket -> sdram_s1_translator_avalon_universal_slave_0_agent:cp_startofpacket
	wire  [107:0] burst_adapter_008_source0_data;                                                                      // burst_adapter_008:source0_data -> sdram_s1_translator_avalon_universal_slave_0_agent:cp_data
	wire          burst_adapter_008_source0_ready;                                                                     // sdram_s1_translator_avalon_universal_slave_0_agent:cp_ready -> burst_adapter_008:source0_ready
	wire    [2:0] burst_adapter_008_source0_channel;                                                                   // burst_adapter_008:source0_channel -> sdram_s1_translator_avalon_universal_slave_0_agent:cp_channel
	wire          width_adapter_cmd_source_endofpacket;                                                                // width_adapter:cmd_out_endofpacket -> hps_0_f2h_axi_slave_agent:write_cp_endofpacket
	wire          width_adapter_cmd_source_valid;                                                                      // width_adapter:cmd_out_valid -> hps_0_f2h_axi_slave_agent:write_cp_valid
	wire          width_adapter_cmd_source_startofpacket;                                                              // width_adapter:cmd_out_startofpacket -> hps_0_f2h_axi_slave_agent:write_cp_startofpacket
	wire  [150:0] width_adapter_cmd_source_data;                                                                       // width_adapter:cmd_out_data -> hps_0_f2h_axi_slave_agent:write_cp_data
	wire    [1:0] width_adapter_cmd_source_channel;                                                                    // width_adapter:cmd_out_channel -> hps_0_f2h_axi_slave_agent:write_cp_channel
	wire          width_adapter_cmd_source_ready;                                                                      // hps_0_f2h_axi_slave_agent:write_cp_ready -> width_adapter:cmd_out_ready
	wire          id_router_src_endofpacket;                                                                           // id_router:src_endofpacket -> width_adapter:rsp_in_endofpacket
	wire          id_router_src_valid;                                                                                 // id_router:src_valid -> width_adapter:rsp_in_valid
	wire          id_router_src_startofpacket;                                                                         // id_router:src_startofpacket -> width_adapter:rsp_in_startofpacket
	wire  [150:0] id_router_src_data;                                                                                  // id_router:src_data -> width_adapter:rsp_in_data
	wire    [1:0] id_router_src_channel;                                                                               // id_router:src_channel -> width_adapter:rsp_in_channel
	wire          id_router_src_ready;                                                                                 // width_adapter:rsp_in_ready -> id_router:src_ready
	wire          width_adapter_001_cmd_source_endofpacket;                                                            // width_adapter_001:cmd_out_endofpacket -> hps_0_f2h_axi_slave_agent:read_cp_endofpacket
	wire          width_adapter_001_cmd_source_valid;                                                                  // width_adapter_001:cmd_out_valid -> hps_0_f2h_axi_slave_agent:read_cp_valid
	wire          width_adapter_001_cmd_source_startofpacket;                                                          // width_adapter_001:cmd_out_startofpacket -> hps_0_f2h_axi_slave_agent:read_cp_startofpacket
	wire  [150:0] width_adapter_001_cmd_source_data;                                                                   // width_adapter_001:cmd_out_data -> hps_0_f2h_axi_slave_agent:read_cp_data
	wire    [1:0] width_adapter_001_cmd_source_channel;                                                                // width_adapter_001:cmd_out_channel -> hps_0_f2h_axi_slave_agent:read_cp_channel
	wire          width_adapter_001_cmd_source_ready;                                                                  // hps_0_f2h_axi_slave_agent:read_cp_ready -> width_adapter_001:cmd_out_ready
	wire          id_router_001_src_endofpacket;                                                                       // id_router_001:src_endofpacket -> width_adapter_001:rsp_in_endofpacket
	wire          id_router_001_src_valid;                                                                             // id_router_001:src_valid -> width_adapter_001:rsp_in_valid
	wire          id_router_001_src_startofpacket;                                                                     // id_router_001:src_startofpacket -> width_adapter_001:rsp_in_startofpacket
	wire  [150:0] id_router_001_src_data;                                                                              // id_router_001:src_data -> width_adapter_001:rsp_in_data
	wire    [1:0] id_router_001_src_channel;                                                                           // id_router_001:src_channel -> width_adapter_001:rsp_in_channel
	wire          id_router_001_src_ready;                                                                             // width_adapter_001:rsp_in_ready -> id_router_001:src_ready
	wire          addr_router_005_src_endofpacket;                                                                     // addr_router_005:src_endofpacket -> width_adapter_002:cmd_in_endofpacket
	wire          addr_router_005_src_valid;                                                                           // addr_router_005:src_valid -> width_adapter_002:cmd_in_valid
	wire          addr_router_005_src_startofpacket;                                                                   // addr_router_005:src_startofpacket -> width_adapter_002:cmd_in_startofpacket
	wire  [125:0] addr_router_005_src_data;                                                                            // addr_router_005:src_data -> width_adapter_002:cmd_in_data
	wire    [2:0] addr_router_005_src_channel;                                                                         // addr_router_005:src_channel -> width_adapter_002:cmd_in_channel
	wire          addr_router_005_src_ready;                                                                           // width_adapter_002:cmd_in_ready -> addr_router_005:src_ready
	wire          width_adapter_002_rsp_source_endofpacket;                                                            // width_adapter_002:rsp_out_endofpacket -> alt_vip_vfr_0_avalon_master_translator_avalon_universal_master_0_agent:rp_endofpacket
	wire          width_adapter_002_rsp_source_valid;                                                                  // width_adapter_002:rsp_out_valid -> alt_vip_vfr_0_avalon_master_translator_avalon_universal_master_0_agent:rp_valid
	wire          width_adapter_002_rsp_source_startofpacket;                                                          // width_adapter_002:rsp_out_startofpacket -> alt_vip_vfr_0_avalon_master_translator_avalon_universal_master_0_agent:rp_startofpacket
	wire  [125:0] width_adapter_002_rsp_source_data;                                                                   // width_adapter_002:rsp_out_data -> alt_vip_vfr_0_avalon_master_translator_avalon_universal_master_0_agent:rp_data
	wire    [2:0] width_adapter_002_rsp_source_channel;                                                                // width_adapter_002:rsp_out_channel -> alt_vip_vfr_0_avalon_master_translator_avalon_universal_master_0_agent:rp_channel
	wire          width_adapter_002_rsp_source_ready;                                                                  // alt_vip_vfr_0_avalon_master_translator_avalon_universal_master_0_agent:rp_ready -> width_adapter_002:rsp_out_ready
	wire          width_adapter_003_cmd_source_endofpacket;                                                            // width_adapter_003:cmd_out_endofpacket -> burst_adapter_008:sink0_endofpacket
	wire          width_adapter_003_cmd_source_valid;                                                                  // width_adapter_003:cmd_out_valid -> burst_adapter_008:sink0_valid
	wire          width_adapter_003_cmd_source_startofpacket;                                                          // width_adapter_003:cmd_out_startofpacket -> burst_adapter_008:sink0_startofpacket
	wire  [107:0] width_adapter_003_cmd_source_data;                                                                   // width_adapter_003:cmd_out_data -> burst_adapter_008:sink0_data
	wire    [2:0] width_adapter_003_cmd_source_channel;                                                                // width_adapter_003:cmd_out_channel -> burst_adapter_008:sink0_channel
	wire          width_adapter_003_cmd_source_ready;                                                                  // burst_adapter_008:sink0_ready -> width_adapter_003:cmd_out_ready
	wire          id_router_010_src_endofpacket;                                                                       // id_router_010:src_endofpacket -> width_adapter_003:rsp_in_endofpacket
	wire          id_router_010_src_valid;                                                                             // id_router_010:src_valid -> width_adapter_003:rsp_in_valid
	wire          id_router_010_src_startofpacket;                                                                     // id_router_010:src_startofpacket -> width_adapter_003:rsp_in_startofpacket
	wire  [107:0] id_router_010_src_data;                                                                              // id_router_010:src_data -> width_adapter_003:rsp_in_data
	wire    [2:0] id_router_010_src_channel;                                                                           // id_router_010:src_channel -> width_adapter_003:rsp_in_channel
	wire          id_router_010_src_ready;                                                                             // width_adapter_003:rsp_in_ready -> id_router_010:src_ready
	wire          rst_controller_reset_out_reset;                                                                      // rst_controller:reset_out -> [addr_router:reset, burst_adapter:reset, burst_adapter_001:reset, burst_adapter_002:reset, burst_adapter_003:reset, burst_adapter_004:reset, button_pio:reset_n, button_pio_s1_translator:reset, button_pio_s1_translator_avalon_universal_slave_0_agent:reset, button_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, cmd_xbar_demux:reset, cmd_xbar_mux_002:reset, cmd_xbar_mux_003:reset, cmd_xbar_mux_004:reset, cmd_xbar_mux_005:reset, cmd_xbar_mux_006:reset, dipsw_pio:reset_n, dipsw_pio_s1_translator:reset, dipsw_pio_s1_translator_avalon_universal_slave_0_agent:reset, dipsw_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, dipsw_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, id_router_002:reset, id_router_003:reset, id_router_004:reset, id_router_005:reset, id_router_006:reset, jtag_uart:rst_n, jtag_uart_avalon_jtag_slave_translator:reset, jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent:reset, jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, led_pio:reset_n, led_pio_s1_translator:reset, led_pio_s1_translator_avalon_universal_slave_0_agent:reset, led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, limiter:reset, master_secure_master_translator:reset, master_secure_master_translator_avalon_universal_master_0_agent:reset, oc_i2c_master_0:wb_rst_i, oc_i2c_master_0_avalon_slave_0_translator:reset, oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent:reset, oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, pll_audio:rst, pll_sdram:rst, pll_stream:rst, rsp_xbar_demux_002:reset, rsp_xbar_demux_003:reset, rsp_xbar_demux_004:reset, rsp_xbar_demux_005:reset, rsp_xbar_demux_006:reset, rsp_xbar_mux:reset]
	wire          rst_controller_001_reset_out_reset;                                                                  // rst_controller_001:reset_out -> [addr_router_005:reset, alt_vip_vfr_0:master_reset, alt_vip_vfr_0_avalon_master_translator:reset, alt_vip_vfr_0_avalon_master_translator_avalon_universal_master_0_agent:reset, burst_adapter_008:reset, cmd_xbar_demux_005:reset, cmd_xbar_mux_010:reset, id_router_010:reset, rsp_xbar_demux_010:reset, sdram:reset_n, sdram_s1_translator:reset, sdram_s1_translator_avalon_universal_slave_0_agent:reset, sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, width_adapter_002:reset, width_adapter_003:reset]
	wire          rst_controller_002_reset_out_reset;                                                                  // rst_controller_002:reset_out -> [LOG_Generate_0:reset, alt_vip_itc_0:rst, alt_vip_mix_0:reset, alt_vip_mix_0_control_translator:reset, alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent:reset, alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, alt_vip_tpg_0:reset, alt_vip_vfr_0:reset, alt_vip_vfr_0_avalon_slave_translator:reset, alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent:reset, alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, avalon_st_adapter:in_rst_0_reset, burst_adapter_005:reset, burst_adapter_006:reset, cmd_xbar_mux_007:reset, cmd_xbar_mux_008:reset, crosser:out_reset, crosser_001:out_reset, crosser_003:out_reset, crosser_004:out_reset, crosser_006:in_reset, crosser_007:in_reset, crosser_008:in_reset, crosser_009:in_reset, id_router_007:reset, id_router_008:reset, rsp_xbar_demux_007:reset, rsp_xbar_demux_008:reset, timing_adapter_0:reset_n]
	wire          rst_controller_003_reset_out_reset;                                                                  // rst_controller_003:reset_out -> [AUDIO_IF_0:avs_s1_reset, AUDIO_IF_0_avalon_slave_translator:reset, AUDIO_IF_0_avalon_slave_translator_avalon_universal_slave_0_agent:reset, AUDIO_IF_0_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo:reset, AUDIO_IF_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo:reset, burst_adapter_007:reset, cmd_xbar_mux_009:reset, crosser_002:out_reset, crosser_005:out_reset, crosser_010:in_reset, crosser_011:in_reset, id_router_009:reset, rsp_xbar_demux_009:reset]
	wire          rst_controller_004_reset_out_reset;                                                                  // rst_controller_004:reset_out -> [addr_router_001:reset, addr_router_002:reset, cmd_xbar_demux_001:reset, cmd_xbar_demux_002:reset, crosser:in_reset, crosser_001:in_reset, crosser_002:in_reset, crosser_003:in_reset, crosser_004:in_reset, crosser_005:in_reset, crosser_006:out_reset, crosser_007:out_reset, crosser_008:out_reset, crosser_009:out_reset, crosser_010:out_reset, crosser_011:out_reset, hps_0_f2h_axi_slave_agent:aresetn, hps_0_h2f_lw_axi_master_agent:aresetn, id_router:reset, id_router_001:reset, limiter_001:reset, limiter_002:reset, rsp_xbar_demux:reset, rsp_xbar_demux_001:reset, rsp_xbar_mux_001:reset, rsp_xbar_mux_002:reset, width_adapter:reset, width_adapter_001:reset]
	wire          rst_controller_005_reset_out_reset;                                                                  // rst_controller_005:reset_out -> [addr_router_003:reset, addr_router_004:reset, cmd_xbar_demux_003:reset, cmd_xbar_demux_004:reset, hps_0_h2f_axi_master_agent:aresetn]
	wire          cmd_xbar_demux_src0_endofpacket;                                                                     // cmd_xbar_demux:src0_endofpacket -> width_adapter:cmd_in_endofpacket
	wire          cmd_xbar_demux_src0_valid;                                                                           // cmd_xbar_demux:src0_valid -> width_adapter:cmd_in_valid
	wire          cmd_xbar_demux_src0_startofpacket;                                                                   // cmd_xbar_demux:src0_startofpacket -> width_adapter:cmd_in_startofpacket
	wire  [114:0] cmd_xbar_demux_src0_data;                                                                            // cmd_xbar_demux:src0_data -> width_adapter:cmd_in_data
	wire    [1:0] cmd_xbar_demux_src0_channel;                                                                         // cmd_xbar_demux:src0_channel -> width_adapter:cmd_in_channel
	wire          cmd_xbar_demux_src1_endofpacket;                                                                     // cmd_xbar_demux:src1_endofpacket -> width_adapter_001:cmd_in_endofpacket
	wire          cmd_xbar_demux_src1_valid;                                                                           // cmd_xbar_demux:src1_valid -> width_adapter_001:cmd_in_valid
	wire          cmd_xbar_demux_src1_startofpacket;                                                                   // cmd_xbar_demux:src1_startofpacket -> width_adapter_001:cmd_in_startofpacket
	wire  [114:0] cmd_xbar_demux_src1_data;                                                                            // cmd_xbar_demux:src1_data -> width_adapter_001:cmd_in_data
	wire    [1:0] cmd_xbar_demux_src1_channel;                                                                         // cmd_xbar_demux:src1_channel -> width_adapter_001:cmd_in_channel
	wire          rsp_xbar_demux_src0_endofpacket;                                                                     // rsp_xbar_demux:src0_endofpacket -> rsp_xbar_mux:sink0_endofpacket
	wire          rsp_xbar_demux_src0_valid;                                                                           // rsp_xbar_demux:src0_valid -> rsp_xbar_mux:sink0_valid
	wire          rsp_xbar_demux_src0_startofpacket;                                                                   // rsp_xbar_demux:src0_startofpacket -> rsp_xbar_mux:sink0_startofpacket
	wire  [114:0] rsp_xbar_demux_src0_data;                                                                            // rsp_xbar_demux:src0_data -> rsp_xbar_mux:sink0_data
	wire    [1:0] rsp_xbar_demux_src0_channel;                                                                         // rsp_xbar_demux:src0_channel -> rsp_xbar_mux:sink0_channel
	wire          rsp_xbar_demux_src0_ready;                                                                           // rsp_xbar_mux:sink0_ready -> rsp_xbar_demux:src0_ready
	wire          rsp_xbar_demux_001_src0_endofpacket;                                                                 // rsp_xbar_demux_001:src0_endofpacket -> rsp_xbar_mux:sink1_endofpacket
	wire          rsp_xbar_demux_001_src0_valid;                                                                       // rsp_xbar_demux_001:src0_valid -> rsp_xbar_mux:sink1_valid
	wire          rsp_xbar_demux_001_src0_startofpacket;                                                               // rsp_xbar_demux_001:src0_startofpacket -> rsp_xbar_mux:sink1_startofpacket
	wire  [114:0] rsp_xbar_demux_001_src0_data;                                                                        // rsp_xbar_demux_001:src0_data -> rsp_xbar_mux:sink1_data
	wire    [1:0] rsp_xbar_demux_001_src0_channel;                                                                     // rsp_xbar_demux_001:src0_channel -> rsp_xbar_mux:sink1_channel
	wire          rsp_xbar_demux_001_src0_ready;                                                                       // rsp_xbar_mux:sink1_ready -> rsp_xbar_demux_001:src0_ready
	wire          limiter_cmd_src_endofpacket;                                                                         // limiter:cmd_src_endofpacket -> cmd_xbar_demux:sink_endofpacket
	wire          limiter_cmd_src_startofpacket;                                                                       // limiter:cmd_src_startofpacket -> cmd_xbar_demux:sink_startofpacket
	wire  [114:0] limiter_cmd_src_data;                                                                                // limiter:cmd_src_data -> cmd_xbar_demux:sink_data
	wire    [1:0] limiter_cmd_src_channel;                                                                             // limiter:cmd_src_channel -> cmd_xbar_demux:sink_channel
	wire          limiter_cmd_src_ready;                                                                               // cmd_xbar_demux:sink_ready -> limiter:cmd_src_ready
	wire          rsp_xbar_mux_src_endofpacket;                                                                        // rsp_xbar_mux:src_endofpacket -> limiter:rsp_sink_endofpacket
	wire          rsp_xbar_mux_src_valid;                                                                              // rsp_xbar_mux:src_valid -> limiter:rsp_sink_valid
	wire          rsp_xbar_mux_src_startofpacket;                                                                      // rsp_xbar_mux:src_startofpacket -> limiter:rsp_sink_startofpacket
	wire  [114:0] rsp_xbar_mux_src_data;                                                                               // rsp_xbar_mux:src_data -> limiter:rsp_sink_data
	wire    [1:0] rsp_xbar_mux_src_channel;                                                                            // rsp_xbar_mux:src_channel -> limiter:rsp_sink_channel
	wire          rsp_xbar_mux_src_ready;                                                                              // limiter:rsp_sink_ready -> rsp_xbar_mux:src_ready
	wire          cmd_xbar_demux_src0_ready;                                                                           // width_adapter:cmd_in_ready -> cmd_xbar_demux:src0_ready
	wire          width_adapter_rsp_source_endofpacket;                                                                // width_adapter:rsp_out_endofpacket -> rsp_xbar_demux:sink_endofpacket
	wire          width_adapter_rsp_source_valid;                                                                      // width_adapter:rsp_out_valid -> rsp_xbar_demux:sink_valid
	wire          width_adapter_rsp_source_startofpacket;                                                              // width_adapter:rsp_out_startofpacket -> rsp_xbar_demux:sink_startofpacket
	wire  [114:0] width_adapter_rsp_source_data;                                                                       // width_adapter:rsp_out_data -> rsp_xbar_demux:sink_data
	wire    [1:0] width_adapter_rsp_source_channel;                                                                    // width_adapter:rsp_out_channel -> rsp_xbar_demux:sink_channel
	wire          width_adapter_rsp_source_ready;                                                                      // rsp_xbar_demux:sink_ready -> width_adapter:rsp_out_ready
	wire          cmd_xbar_demux_src1_ready;                                                                           // width_adapter_001:cmd_in_ready -> cmd_xbar_demux:src1_ready
	wire          width_adapter_001_rsp_source_endofpacket;                                                            // width_adapter_001:rsp_out_endofpacket -> rsp_xbar_demux_001:sink_endofpacket
	wire          width_adapter_001_rsp_source_valid;                                                                  // width_adapter_001:rsp_out_valid -> rsp_xbar_demux_001:sink_valid
	wire          width_adapter_001_rsp_source_startofpacket;                                                          // width_adapter_001:rsp_out_startofpacket -> rsp_xbar_demux_001:sink_startofpacket
	wire  [114:0] width_adapter_001_rsp_source_data;                                                                   // width_adapter_001:rsp_out_data -> rsp_xbar_demux_001:sink_data
	wire    [1:0] width_adapter_001_rsp_source_channel;                                                                // width_adapter_001:rsp_out_channel -> rsp_xbar_demux_001:sink_channel
	wire          width_adapter_001_rsp_source_ready;                                                                  // rsp_xbar_demux_001:sink_ready -> width_adapter_001:rsp_out_ready
	wire          cmd_xbar_demux_001_src0_endofpacket;                                                                 // cmd_xbar_demux_001:src0_endofpacket -> cmd_xbar_mux_002:sink0_endofpacket
	wire          cmd_xbar_demux_001_src0_valid;                                                                       // cmd_xbar_demux_001:src0_valid -> cmd_xbar_mux_002:sink0_valid
	wire          cmd_xbar_demux_001_src0_startofpacket;                                                               // cmd_xbar_demux_001:src0_startofpacket -> cmd_xbar_mux_002:sink0_startofpacket
	wire  [112:0] cmd_xbar_demux_001_src0_data;                                                                        // cmd_xbar_demux_001:src0_data -> cmd_xbar_mux_002:sink0_data
	wire    [7:0] cmd_xbar_demux_001_src0_channel;                                                                     // cmd_xbar_demux_001:src0_channel -> cmd_xbar_mux_002:sink0_channel
	wire          cmd_xbar_demux_001_src0_ready;                                                                       // cmd_xbar_mux_002:sink0_ready -> cmd_xbar_demux_001:src0_ready
	wire          cmd_xbar_demux_001_src1_endofpacket;                                                                 // cmd_xbar_demux_001:src1_endofpacket -> cmd_xbar_mux_003:sink0_endofpacket
	wire          cmd_xbar_demux_001_src1_valid;                                                                       // cmd_xbar_demux_001:src1_valid -> cmd_xbar_mux_003:sink0_valid
	wire          cmd_xbar_demux_001_src1_startofpacket;                                                               // cmd_xbar_demux_001:src1_startofpacket -> cmd_xbar_mux_003:sink0_startofpacket
	wire  [112:0] cmd_xbar_demux_001_src1_data;                                                                        // cmd_xbar_demux_001:src1_data -> cmd_xbar_mux_003:sink0_data
	wire    [7:0] cmd_xbar_demux_001_src1_channel;                                                                     // cmd_xbar_demux_001:src1_channel -> cmd_xbar_mux_003:sink0_channel
	wire          cmd_xbar_demux_001_src1_ready;                                                                       // cmd_xbar_mux_003:sink0_ready -> cmd_xbar_demux_001:src1_ready
	wire          cmd_xbar_demux_001_src2_endofpacket;                                                                 // cmd_xbar_demux_001:src2_endofpacket -> cmd_xbar_mux_004:sink0_endofpacket
	wire          cmd_xbar_demux_001_src2_valid;                                                                       // cmd_xbar_demux_001:src2_valid -> cmd_xbar_mux_004:sink0_valid
	wire          cmd_xbar_demux_001_src2_startofpacket;                                                               // cmd_xbar_demux_001:src2_startofpacket -> cmd_xbar_mux_004:sink0_startofpacket
	wire  [112:0] cmd_xbar_demux_001_src2_data;                                                                        // cmd_xbar_demux_001:src2_data -> cmd_xbar_mux_004:sink0_data
	wire    [7:0] cmd_xbar_demux_001_src2_channel;                                                                     // cmd_xbar_demux_001:src2_channel -> cmd_xbar_mux_004:sink0_channel
	wire          cmd_xbar_demux_001_src2_ready;                                                                       // cmd_xbar_mux_004:sink0_ready -> cmd_xbar_demux_001:src2_ready
	wire          cmd_xbar_demux_001_src3_endofpacket;                                                                 // cmd_xbar_demux_001:src3_endofpacket -> cmd_xbar_mux_005:sink0_endofpacket
	wire          cmd_xbar_demux_001_src3_valid;                                                                       // cmd_xbar_demux_001:src3_valid -> cmd_xbar_mux_005:sink0_valid
	wire          cmd_xbar_demux_001_src3_startofpacket;                                                               // cmd_xbar_demux_001:src3_startofpacket -> cmd_xbar_mux_005:sink0_startofpacket
	wire  [112:0] cmd_xbar_demux_001_src3_data;                                                                        // cmd_xbar_demux_001:src3_data -> cmd_xbar_mux_005:sink0_data
	wire    [7:0] cmd_xbar_demux_001_src3_channel;                                                                     // cmd_xbar_demux_001:src3_channel -> cmd_xbar_mux_005:sink0_channel
	wire          cmd_xbar_demux_001_src3_ready;                                                                       // cmd_xbar_mux_005:sink0_ready -> cmd_xbar_demux_001:src3_ready
	wire          cmd_xbar_demux_001_src4_endofpacket;                                                                 // cmd_xbar_demux_001:src4_endofpacket -> cmd_xbar_mux_006:sink0_endofpacket
	wire          cmd_xbar_demux_001_src4_valid;                                                                       // cmd_xbar_demux_001:src4_valid -> cmd_xbar_mux_006:sink0_valid
	wire          cmd_xbar_demux_001_src4_startofpacket;                                                               // cmd_xbar_demux_001:src4_startofpacket -> cmd_xbar_mux_006:sink0_startofpacket
	wire  [112:0] cmd_xbar_demux_001_src4_data;                                                                        // cmd_xbar_demux_001:src4_data -> cmd_xbar_mux_006:sink0_data
	wire    [7:0] cmd_xbar_demux_001_src4_channel;                                                                     // cmd_xbar_demux_001:src4_channel -> cmd_xbar_mux_006:sink0_channel
	wire          cmd_xbar_demux_001_src4_ready;                                                                       // cmd_xbar_mux_006:sink0_ready -> cmd_xbar_demux_001:src4_ready
	wire          cmd_xbar_demux_002_src0_endofpacket;                                                                 // cmd_xbar_demux_002:src0_endofpacket -> cmd_xbar_mux_002:sink1_endofpacket
	wire          cmd_xbar_demux_002_src0_valid;                                                                       // cmd_xbar_demux_002:src0_valid -> cmd_xbar_mux_002:sink1_valid
	wire          cmd_xbar_demux_002_src0_startofpacket;                                                               // cmd_xbar_demux_002:src0_startofpacket -> cmd_xbar_mux_002:sink1_startofpacket
	wire  [112:0] cmd_xbar_demux_002_src0_data;                                                                        // cmd_xbar_demux_002:src0_data -> cmd_xbar_mux_002:sink1_data
	wire    [7:0] cmd_xbar_demux_002_src0_channel;                                                                     // cmd_xbar_demux_002:src0_channel -> cmd_xbar_mux_002:sink1_channel
	wire          cmd_xbar_demux_002_src0_ready;                                                                       // cmd_xbar_mux_002:sink1_ready -> cmd_xbar_demux_002:src0_ready
	wire          cmd_xbar_demux_002_src1_endofpacket;                                                                 // cmd_xbar_demux_002:src1_endofpacket -> cmd_xbar_mux_003:sink1_endofpacket
	wire          cmd_xbar_demux_002_src1_valid;                                                                       // cmd_xbar_demux_002:src1_valid -> cmd_xbar_mux_003:sink1_valid
	wire          cmd_xbar_demux_002_src1_startofpacket;                                                               // cmd_xbar_demux_002:src1_startofpacket -> cmd_xbar_mux_003:sink1_startofpacket
	wire  [112:0] cmd_xbar_demux_002_src1_data;                                                                        // cmd_xbar_demux_002:src1_data -> cmd_xbar_mux_003:sink1_data
	wire    [7:0] cmd_xbar_demux_002_src1_channel;                                                                     // cmd_xbar_demux_002:src1_channel -> cmd_xbar_mux_003:sink1_channel
	wire          cmd_xbar_demux_002_src1_ready;                                                                       // cmd_xbar_mux_003:sink1_ready -> cmd_xbar_demux_002:src1_ready
	wire          cmd_xbar_demux_002_src2_endofpacket;                                                                 // cmd_xbar_demux_002:src2_endofpacket -> cmd_xbar_mux_004:sink1_endofpacket
	wire          cmd_xbar_demux_002_src2_valid;                                                                       // cmd_xbar_demux_002:src2_valid -> cmd_xbar_mux_004:sink1_valid
	wire          cmd_xbar_demux_002_src2_startofpacket;                                                               // cmd_xbar_demux_002:src2_startofpacket -> cmd_xbar_mux_004:sink1_startofpacket
	wire  [112:0] cmd_xbar_demux_002_src2_data;                                                                        // cmd_xbar_demux_002:src2_data -> cmd_xbar_mux_004:sink1_data
	wire    [7:0] cmd_xbar_demux_002_src2_channel;                                                                     // cmd_xbar_demux_002:src2_channel -> cmd_xbar_mux_004:sink1_channel
	wire          cmd_xbar_demux_002_src2_ready;                                                                       // cmd_xbar_mux_004:sink1_ready -> cmd_xbar_demux_002:src2_ready
	wire          cmd_xbar_demux_002_src3_endofpacket;                                                                 // cmd_xbar_demux_002:src3_endofpacket -> cmd_xbar_mux_005:sink1_endofpacket
	wire          cmd_xbar_demux_002_src3_valid;                                                                       // cmd_xbar_demux_002:src3_valid -> cmd_xbar_mux_005:sink1_valid
	wire          cmd_xbar_demux_002_src3_startofpacket;                                                               // cmd_xbar_demux_002:src3_startofpacket -> cmd_xbar_mux_005:sink1_startofpacket
	wire  [112:0] cmd_xbar_demux_002_src3_data;                                                                        // cmd_xbar_demux_002:src3_data -> cmd_xbar_mux_005:sink1_data
	wire    [7:0] cmd_xbar_demux_002_src3_channel;                                                                     // cmd_xbar_demux_002:src3_channel -> cmd_xbar_mux_005:sink1_channel
	wire          cmd_xbar_demux_002_src3_ready;                                                                       // cmd_xbar_mux_005:sink1_ready -> cmd_xbar_demux_002:src3_ready
	wire          cmd_xbar_demux_002_src4_endofpacket;                                                                 // cmd_xbar_demux_002:src4_endofpacket -> cmd_xbar_mux_006:sink1_endofpacket
	wire          cmd_xbar_demux_002_src4_valid;                                                                       // cmd_xbar_demux_002:src4_valid -> cmd_xbar_mux_006:sink1_valid
	wire          cmd_xbar_demux_002_src4_startofpacket;                                                               // cmd_xbar_demux_002:src4_startofpacket -> cmd_xbar_mux_006:sink1_startofpacket
	wire  [112:0] cmd_xbar_demux_002_src4_data;                                                                        // cmd_xbar_demux_002:src4_data -> cmd_xbar_mux_006:sink1_data
	wire    [7:0] cmd_xbar_demux_002_src4_channel;                                                                     // cmd_xbar_demux_002:src4_channel -> cmd_xbar_mux_006:sink1_channel
	wire          cmd_xbar_demux_002_src4_ready;                                                                       // cmd_xbar_mux_006:sink1_ready -> cmd_xbar_demux_002:src4_ready
	wire          rsp_xbar_demux_002_src0_endofpacket;                                                                 // rsp_xbar_demux_002:src0_endofpacket -> rsp_xbar_mux_001:sink0_endofpacket
	wire          rsp_xbar_demux_002_src0_valid;                                                                       // rsp_xbar_demux_002:src0_valid -> rsp_xbar_mux_001:sink0_valid
	wire          rsp_xbar_demux_002_src0_startofpacket;                                                               // rsp_xbar_demux_002:src0_startofpacket -> rsp_xbar_mux_001:sink0_startofpacket
	wire  [112:0] rsp_xbar_demux_002_src0_data;                                                                        // rsp_xbar_demux_002:src0_data -> rsp_xbar_mux_001:sink0_data
	wire    [7:0] rsp_xbar_demux_002_src0_channel;                                                                     // rsp_xbar_demux_002:src0_channel -> rsp_xbar_mux_001:sink0_channel
	wire          rsp_xbar_demux_002_src0_ready;                                                                       // rsp_xbar_mux_001:sink0_ready -> rsp_xbar_demux_002:src0_ready
	wire          rsp_xbar_demux_002_src1_endofpacket;                                                                 // rsp_xbar_demux_002:src1_endofpacket -> rsp_xbar_mux_002:sink0_endofpacket
	wire          rsp_xbar_demux_002_src1_valid;                                                                       // rsp_xbar_demux_002:src1_valid -> rsp_xbar_mux_002:sink0_valid
	wire          rsp_xbar_demux_002_src1_startofpacket;                                                               // rsp_xbar_demux_002:src1_startofpacket -> rsp_xbar_mux_002:sink0_startofpacket
	wire  [112:0] rsp_xbar_demux_002_src1_data;                                                                        // rsp_xbar_demux_002:src1_data -> rsp_xbar_mux_002:sink0_data
	wire    [7:0] rsp_xbar_demux_002_src1_channel;                                                                     // rsp_xbar_demux_002:src1_channel -> rsp_xbar_mux_002:sink0_channel
	wire          rsp_xbar_demux_002_src1_ready;                                                                       // rsp_xbar_mux_002:sink0_ready -> rsp_xbar_demux_002:src1_ready
	wire          rsp_xbar_demux_003_src0_endofpacket;                                                                 // rsp_xbar_demux_003:src0_endofpacket -> rsp_xbar_mux_001:sink1_endofpacket
	wire          rsp_xbar_demux_003_src0_valid;                                                                       // rsp_xbar_demux_003:src0_valid -> rsp_xbar_mux_001:sink1_valid
	wire          rsp_xbar_demux_003_src0_startofpacket;                                                               // rsp_xbar_demux_003:src0_startofpacket -> rsp_xbar_mux_001:sink1_startofpacket
	wire  [112:0] rsp_xbar_demux_003_src0_data;                                                                        // rsp_xbar_demux_003:src0_data -> rsp_xbar_mux_001:sink1_data
	wire    [7:0] rsp_xbar_demux_003_src0_channel;                                                                     // rsp_xbar_demux_003:src0_channel -> rsp_xbar_mux_001:sink1_channel
	wire          rsp_xbar_demux_003_src0_ready;                                                                       // rsp_xbar_mux_001:sink1_ready -> rsp_xbar_demux_003:src0_ready
	wire          rsp_xbar_demux_003_src1_endofpacket;                                                                 // rsp_xbar_demux_003:src1_endofpacket -> rsp_xbar_mux_002:sink1_endofpacket
	wire          rsp_xbar_demux_003_src1_valid;                                                                       // rsp_xbar_demux_003:src1_valid -> rsp_xbar_mux_002:sink1_valid
	wire          rsp_xbar_demux_003_src1_startofpacket;                                                               // rsp_xbar_demux_003:src1_startofpacket -> rsp_xbar_mux_002:sink1_startofpacket
	wire  [112:0] rsp_xbar_demux_003_src1_data;                                                                        // rsp_xbar_demux_003:src1_data -> rsp_xbar_mux_002:sink1_data
	wire    [7:0] rsp_xbar_demux_003_src1_channel;                                                                     // rsp_xbar_demux_003:src1_channel -> rsp_xbar_mux_002:sink1_channel
	wire          rsp_xbar_demux_003_src1_ready;                                                                       // rsp_xbar_mux_002:sink1_ready -> rsp_xbar_demux_003:src1_ready
	wire          rsp_xbar_demux_004_src0_endofpacket;                                                                 // rsp_xbar_demux_004:src0_endofpacket -> rsp_xbar_mux_001:sink2_endofpacket
	wire          rsp_xbar_demux_004_src0_valid;                                                                       // rsp_xbar_demux_004:src0_valid -> rsp_xbar_mux_001:sink2_valid
	wire          rsp_xbar_demux_004_src0_startofpacket;                                                               // rsp_xbar_demux_004:src0_startofpacket -> rsp_xbar_mux_001:sink2_startofpacket
	wire  [112:0] rsp_xbar_demux_004_src0_data;                                                                        // rsp_xbar_demux_004:src0_data -> rsp_xbar_mux_001:sink2_data
	wire    [7:0] rsp_xbar_demux_004_src0_channel;                                                                     // rsp_xbar_demux_004:src0_channel -> rsp_xbar_mux_001:sink2_channel
	wire          rsp_xbar_demux_004_src0_ready;                                                                       // rsp_xbar_mux_001:sink2_ready -> rsp_xbar_demux_004:src0_ready
	wire          rsp_xbar_demux_004_src1_endofpacket;                                                                 // rsp_xbar_demux_004:src1_endofpacket -> rsp_xbar_mux_002:sink2_endofpacket
	wire          rsp_xbar_demux_004_src1_valid;                                                                       // rsp_xbar_demux_004:src1_valid -> rsp_xbar_mux_002:sink2_valid
	wire          rsp_xbar_demux_004_src1_startofpacket;                                                               // rsp_xbar_demux_004:src1_startofpacket -> rsp_xbar_mux_002:sink2_startofpacket
	wire  [112:0] rsp_xbar_demux_004_src1_data;                                                                        // rsp_xbar_demux_004:src1_data -> rsp_xbar_mux_002:sink2_data
	wire    [7:0] rsp_xbar_demux_004_src1_channel;                                                                     // rsp_xbar_demux_004:src1_channel -> rsp_xbar_mux_002:sink2_channel
	wire          rsp_xbar_demux_004_src1_ready;                                                                       // rsp_xbar_mux_002:sink2_ready -> rsp_xbar_demux_004:src1_ready
	wire          rsp_xbar_demux_005_src0_endofpacket;                                                                 // rsp_xbar_demux_005:src0_endofpacket -> rsp_xbar_mux_001:sink3_endofpacket
	wire          rsp_xbar_demux_005_src0_valid;                                                                       // rsp_xbar_demux_005:src0_valid -> rsp_xbar_mux_001:sink3_valid
	wire          rsp_xbar_demux_005_src0_startofpacket;                                                               // rsp_xbar_demux_005:src0_startofpacket -> rsp_xbar_mux_001:sink3_startofpacket
	wire  [112:0] rsp_xbar_demux_005_src0_data;                                                                        // rsp_xbar_demux_005:src0_data -> rsp_xbar_mux_001:sink3_data
	wire    [7:0] rsp_xbar_demux_005_src0_channel;                                                                     // rsp_xbar_demux_005:src0_channel -> rsp_xbar_mux_001:sink3_channel
	wire          rsp_xbar_demux_005_src0_ready;                                                                       // rsp_xbar_mux_001:sink3_ready -> rsp_xbar_demux_005:src0_ready
	wire          rsp_xbar_demux_005_src1_endofpacket;                                                                 // rsp_xbar_demux_005:src1_endofpacket -> rsp_xbar_mux_002:sink3_endofpacket
	wire          rsp_xbar_demux_005_src1_valid;                                                                       // rsp_xbar_demux_005:src1_valid -> rsp_xbar_mux_002:sink3_valid
	wire          rsp_xbar_demux_005_src1_startofpacket;                                                               // rsp_xbar_demux_005:src1_startofpacket -> rsp_xbar_mux_002:sink3_startofpacket
	wire  [112:0] rsp_xbar_demux_005_src1_data;                                                                        // rsp_xbar_demux_005:src1_data -> rsp_xbar_mux_002:sink3_data
	wire    [7:0] rsp_xbar_demux_005_src1_channel;                                                                     // rsp_xbar_demux_005:src1_channel -> rsp_xbar_mux_002:sink3_channel
	wire          rsp_xbar_demux_005_src1_ready;                                                                       // rsp_xbar_mux_002:sink3_ready -> rsp_xbar_demux_005:src1_ready
	wire          rsp_xbar_demux_006_src0_endofpacket;                                                                 // rsp_xbar_demux_006:src0_endofpacket -> rsp_xbar_mux_001:sink4_endofpacket
	wire          rsp_xbar_demux_006_src0_valid;                                                                       // rsp_xbar_demux_006:src0_valid -> rsp_xbar_mux_001:sink4_valid
	wire          rsp_xbar_demux_006_src0_startofpacket;                                                               // rsp_xbar_demux_006:src0_startofpacket -> rsp_xbar_mux_001:sink4_startofpacket
	wire  [112:0] rsp_xbar_demux_006_src0_data;                                                                        // rsp_xbar_demux_006:src0_data -> rsp_xbar_mux_001:sink4_data
	wire    [7:0] rsp_xbar_demux_006_src0_channel;                                                                     // rsp_xbar_demux_006:src0_channel -> rsp_xbar_mux_001:sink4_channel
	wire          rsp_xbar_demux_006_src0_ready;                                                                       // rsp_xbar_mux_001:sink4_ready -> rsp_xbar_demux_006:src0_ready
	wire          rsp_xbar_demux_006_src1_endofpacket;                                                                 // rsp_xbar_demux_006:src1_endofpacket -> rsp_xbar_mux_002:sink4_endofpacket
	wire          rsp_xbar_demux_006_src1_valid;                                                                       // rsp_xbar_demux_006:src1_valid -> rsp_xbar_mux_002:sink4_valid
	wire          rsp_xbar_demux_006_src1_startofpacket;                                                               // rsp_xbar_demux_006:src1_startofpacket -> rsp_xbar_mux_002:sink4_startofpacket
	wire  [112:0] rsp_xbar_demux_006_src1_data;                                                                        // rsp_xbar_demux_006:src1_data -> rsp_xbar_mux_002:sink4_data
	wire    [7:0] rsp_xbar_demux_006_src1_channel;                                                                     // rsp_xbar_demux_006:src1_channel -> rsp_xbar_mux_002:sink4_channel
	wire          rsp_xbar_demux_006_src1_ready;                                                                       // rsp_xbar_mux_002:sink4_ready -> rsp_xbar_demux_006:src1_ready
	wire          limiter_001_cmd_src_endofpacket;                                                                     // limiter_001:cmd_src_endofpacket -> cmd_xbar_demux_001:sink_endofpacket
	wire          limiter_001_cmd_src_startofpacket;                                                                   // limiter_001:cmd_src_startofpacket -> cmd_xbar_demux_001:sink_startofpacket
	wire  [112:0] limiter_001_cmd_src_data;                                                                            // limiter_001:cmd_src_data -> cmd_xbar_demux_001:sink_data
	wire    [7:0] limiter_001_cmd_src_channel;                                                                         // limiter_001:cmd_src_channel -> cmd_xbar_demux_001:sink_channel
	wire          limiter_001_cmd_src_ready;                                                                           // cmd_xbar_demux_001:sink_ready -> limiter_001:cmd_src_ready
	wire          rsp_xbar_mux_001_src_endofpacket;                                                                    // rsp_xbar_mux_001:src_endofpacket -> limiter_001:rsp_sink_endofpacket
	wire          rsp_xbar_mux_001_src_valid;                                                                          // rsp_xbar_mux_001:src_valid -> limiter_001:rsp_sink_valid
	wire          rsp_xbar_mux_001_src_startofpacket;                                                                  // rsp_xbar_mux_001:src_startofpacket -> limiter_001:rsp_sink_startofpacket
	wire  [112:0] rsp_xbar_mux_001_src_data;                                                                           // rsp_xbar_mux_001:src_data -> limiter_001:rsp_sink_data
	wire    [7:0] rsp_xbar_mux_001_src_channel;                                                                        // rsp_xbar_mux_001:src_channel -> limiter_001:rsp_sink_channel
	wire          rsp_xbar_mux_001_src_ready;                                                                          // limiter_001:rsp_sink_ready -> rsp_xbar_mux_001:src_ready
	wire          limiter_002_cmd_src_endofpacket;                                                                     // limiter_002:cmd_src_endofpacket -> cmd_xbar_demux_002:sink_endofpacket
	wire          limiter_002_cmd_src_startofpacket;                                                                   // limiter_002:cmd_src_startofpacket -> cmd_xbar_demux_002:sink_startofpacket
	wire  [112:0] limiter_002_cmd_src_data;                                                                            // limiter_002:cmd_src_data -> cmd_xbar_demux_002:sink_data
	wire    [7:0] limiter_002_cmd_src_channel;                                                                         // limiter_002:cmd_src_channel -> cmd_xbar_demux_002:sink_channel
	wire          limiter_002_cmd_src_ready;                                                                           // cmd_xbar_demux_002:sink_ready -> limiter_002:cmd_src_ready
	wire          rsp_xbar_mux_002_src_endofpacket;                                                                    // rsp_xbar_mux_002:src_endofpacket -> limiter_002:rsp_sink_endofpacket
	wire          rsp_xbar_mux_002_src_valid;                                                                          // rsp_xbar_mux_002:src_valid -> limiter_002:rsp_sink_valid
	wire          rsp_xbar_mux_002_src_startofpacket;                                                                  // rsp_xbar_mux_002:src_startofpacket -> limiter_002:rsp_sink_startofpacket
	wire  [112:0] rsp_xbar_mux_002_src_data;                                                                           // rsp_xbar_mux_002:src_data -> limiter_002:rsp_sink_data
	wire    [7:0] rsp_xbar_mux_002_src_channel;                                                                        // rsp_xbar_mux_002:src_channel -> limiter_002:rsp_sink_channel
	wire          rsp_xbar_mux_002_src_ready;                                                                          // limiter_002:rsp_sink_ready -> rsp_xbar_mux_002:src_ready
	wire          cmd_xbar_mux_002_src_endofpacket;                                                                    // cmd_xbar_mux_002:src_endofpacket -> burst_adapter:sink0_endofpacket
	wire          cmd_xbar_mux_002_src_valid;                                                                          // cmd_xbar_mux_002:src_valid -> burst_adapter:sink0_valid
	wire          cmd_xbar_mux_002_src_startofpacket;                                                                  // cmd_xbar_mux_002:src_startofpacket -> burst_adapter:sink0_startofpacket
	wire  [112:0] cmd_xbar_mux_002_src_data;                                                                           // cmd_xbar_mux_002:src_data -> burst_adapter:sink0_data
	wire    [7:0] cmd_xbar_mux_002_src_channel;                                                                        // cmd_xbar_mux_002:src_channel -> burst_adapter:sink0_channel
	wire          cmd_xbar_mux_002_src_ready;                                                                          // burst_adapter:sink0_ready -> cmd_xbar_mux_002:src_ready
	wire          id_router_002_src_endofpacket;                                                                       // id_router_002:src_endofpacket -> rsp_xbar_demux_002:sink_endofpacket
	wire          id_router_002_src_valid;                                                                             // id_router_002:src_valid -> rsp_xbar_demux_002:sink_valid
	wire          id_router_002_src_startofpacket;                                                                     // id_router_002:src_startofpacket -> rsp_xbar_demux_002:sink_startofpacket
	wire  [112:0] id_router_002_src_data;                                                                              // id_router_002:src_data -> rsp_xbar_demux_002:sink_data
	wire    [7:0] id_router_002_src_channel;                                                                           // id_router_002:src_channel -> rsp_xbar_demux_002:sink_channel
	wire          id_router_002_src_ready;                                                                             // rsp_xbar_demux_002:sink_ready -> id_router_002:src_ready
	wire          cmd_xbar_mux_003_src_endofpacket;                                                                    // cmd_xbar_mux_003:src_endofpacket -> burst_adapter_001:sink0_endofpacket
	wire          cmd_xbar_mux_003_src_valid;                                                                          // cmd_xbar_mux_003:src_valid -> burst_adapter_001:sink0_valid
	wire          cmd_xbar_mux_003_src_startofpacket;                                                                  // cmd_xbar_mux_003:src_startofpacket -> burst_adapter_001:sink0_startofpacket
	wire  [112:0] cmd_xbar_mux_003_src_data;                                                                           // cmd_xbar_mux_003:src_data -> burst_adapter_001:sink0_data
	wire    [7:0] cmd_xbar_mux_003_src_channel;                                                                        // cmd_xbar_mux_003:src_channel -> burst_adapter_001:sink0_channel
	wire          cmd_xbar_mux_003_src_ready;                                                                          // burst_adapter_001:sink0_ready -> cmd_xbar_mux_003:src_ready
	wire          id_router_003_src_endofpacket;                                                                       // id_router_003:src_endofpacket -> rsp_xbar_demux_003:sink_endofpacket
	wire          id_router_003_src_valid;                                                                             // id_router_003:src_valid -> rsp_xbar_demux_003:sink_valid
	wire          id_router_003_src_startofpacket;                                                                     // id_router_003:src_startofpacket -> rsp_xbar_demux_003:sink_startofpacket
	wire  [112:0] id_router_003_src_data;                                                                              // id_router_003:src_data -> rsp_xbar_demux_003:sink_data
	wire    [7:0] id_router_003_src_channel;                                                                           // id_router_003:src_channel -> rsp_xbar_demux_003:sink_channel
	wire          id_router_003_src_ready;                                                                             // rsp_xbar_demux_003:sink_ready -> id_router_003:src_ready
	wire          cmd_xbar_mux_004_src_endofpacket;                                                                    // cmd_xbar_mux_004:src_endofpacket -> burst_adapter_002:sink0_endofpacket
	wire          cmd_xbar_mux_004_src_valid;                                                                          // cmd_xbar_mux_004:src_valid -> burst_adapter_002:sink0_valid
	wire          cmd_xbar_mux_004_src_startofpacket;                                                                  // cmd_xbar_mux_004:src_startofpacket -> burst_adapter_002:sink0_startofpacket
	wire  [112:0] cmd_xbar_mux_004_src_data;                                                                           // cmd_xbar_mux_004:src_data -> burst_adapter_002:sink0_data
	wire    [7:0] cmd_xbar_mux_004_src_channel;                                                                        // cmd_xbar_mux_004:src_channel -> burst_adapter_002:sink0_channel
	wire          cmd_xbar_mux_004_src_ready;                                                                          // burst_adapter_002:sink0_ready -> cmd_xbar_mux_004:src_ready
	wire          id_router_004_src_endofpacket;                                                                       // id_router_004:src_endofpacket -> rsp_xbar_demux_004:sink_endofpacket
	wire          id_router_004_src_valid;                                                                             // id_router_004:src_valid -> rsp_xbar_demux_004:sink_valid
	wire          id_router_004_src_startofpacket;                                                                     // id_router_004:src_startofpacket -> rsp_xbar_demux_004:sink_startofpacket
	wire  [112:0] id_router_004_src_data;                                                                              // id_router_004:src_data -> rsp_xbar_demux_004:sink_data
	wire    [7:0] id_router_004_src_channel;                                                                           // id_router_004:src_channel -> rsp_xbar_demux_004:sink_channel
	wire          id_router_004_src_ready;                                                                             // rsp_xbar_demux_004:sink_ready -> id_router_004:src_ready
	wire          cmd_xbar_mux_005_src_endofpacket;                                                                    // cmd_xbar_mux_005:src_endofpacket -> burst_adapter_003:sink0_endofpacket
	wire          cmd_xbar_mux_005_src_valid;                                                                          // cmd_xbar_mux_005:src_valid -> burst_adapter_003:sink0_valid
	wire          cmd_xbar_mux_005_src_startofpacket;                                                                  // cmd_xbar_mux_005:src_startofpacket -> burst_adapter_003:sink0_startofpacket
	wire  [112:0] cmd_xbar_mux_005_src_data;                                                                           // cmd_xbar_mux_005:src_data -> burst_adapter_003:sink0_data
	wire    [7:0] cmd_xbar_mux_005_src_channel;                                                                        // cmd_xbar_mux_005:src_channel -> burst_adapter_003:sink0_channel
	wire          cmd_xbar_mux_005_src_ready;                                                                          // burst_adapter_003:sink0_ready -> cmd_xbar_mux_005:src_ready
	wire          id_router_005_src_endofpacket;                                                                       // id_router_005:src_endofpacket -> rsp_xbar_demux_005:sink_endofpacket
	wire          id_router_005_src_valid;                                                                             // id_router_005:src_valid -> rsp_xbar_demux_005:sink_valid
	wire          id_router_005_src_startofpacket;                                                                     // id_router_005:src_startofpacket -> rsp_xbar_demux_005:sink_startofpacket
	wire  [112:0] id_router_005_src_data;                                                                              // id_router_005:src_data -> rsp_xbar_demux_005:sink_data
	wire    [7:0] id_router_005_src_channel;                                                                           // id_router_005:src_channel -> rsp_xbar_demux_005:sink_channel
	wire          id_router_005_src_ready;                                                                             // rsp_xbar_demux_005:sink_ready -> id_router_005:src_ready
	wire          cmd_xbar_mux_006_src_endofpacket;                                                                    // cmd_xbar_mux_006:src_endofpacket -> burst_adapter_004:sink0_endofpacket
	wire          cmd_xbar_mux_006_src_valid;                                                                          // cmd_xbar_mux_006:src_valid -> burst_adapter_004:sink0_valid
	wire          cmd_xbar_mux_006_src_startofpacket;                                                                  // cmd_xbar_mux_006:src_startofpacket -> burst_adapter_004:sink0_startofpacket
	wire  [112:0] cmd_xbar_mux_006_src_data;                                                                           // cmd_xbar_mux_006:src_data -> burst_adapter_004:sink0_data
	wire    [7:0] cmd_xbar_mux_006_src_channel;                                                                        // cmd_xbar_mux_006:src_channel -> burst_adapter_004:sink0_channel
	wire          cmd_xbar_mux_006_src_ready;                                                                          // burst_adapter_004:sink0_ready -> cmd_xbar_mux_006:src_ready
	wire          id_router_006_src_endofpacket;                                                                       // id_router_006:src_endofpacket -> rsp_xbar_demux_006:sink_endofpacket
	wire          id_router_006_src_valid;                                                                             // id_router_006:src_valid -> rsp_xbar_demux_006:sink_valid
	wire          id_router_006_src_startofpacket;                                                                     // id_router_006:src_startofpacket -> rsp_xbar_demux_006:sink_startofpacket
	wire  [112:0] id_router_006_src_data;                                                                              // id_router_006:src_data -> rsp_xbar_demux_006:sink_data
	wire    [7:0] id_router_006_src_channel;                                                                           // id_router_006:src_channel -> rsp_xbar_demux_006:sink_channel
	wire          id_router_006_src_ready;                                                                             // rsp_xbar_demux_006:sink_ready -> id_router_006:src_ready
	wire          cmd_xbar_mux_007_src_endofpacket;                                                                    // cmd_xbar_mux_007:src_endofpacket -> burst_adapter_005:sink0_endofpacket
	wire          cmd_xbar_mux_007_src_valid;                                                                          // cmd_xbar_mux_007:src_valid -> burst_adapter_005:sink0_valid
	wire          cmd_xbar_mux_007_src_startofpacket;                                                                  // cmd_xbar_mux_007:src_startofpacket -> burst_adapter_005:sink0_startofpacket
	wire  [112:0] cmd_xbar_mux_007_src_data;                                                                           // cmd_xbar_mux_007:src_data -> burst_adapter_005:sink0_data
	wire    [7:0] cmd_xbar_mux_007_src_channel;                                                                        // cmd_xbar_mux_007:src_channel -> burst_adapter_005:sink0_channel
	wire          cmd_xbar_mux_007_src_ready;                                                                          // burst_adapter_005:sink0_ready -> cmd_xbar_mux_007:src_ready
	wire          id_router_007_src_endofpacket;                                                                       // id_router_007:src_endofpacket -> rsp_xbar_demux_007:sink_endofpacket
	wire          id_router_007_src_valid;                                                                             // id_router_007:src_valid -> rsp_xbar_demux_007:sink_valid
	wire          id_router_007_src_startofpacket;                                                                     // id_router_007:src_startofpacket -> rsp_xbar_demux_007:sink_startofpacket
	wire  [112:0] id_router_007_src_data;                                                                              // id_router_007:src_data -> rsp_xbar_demux_007:sink_data
	wire    [7:0] id_router_007_src_channel;                                                                           // id_router_007:src_channel -> rsp_xbar_demux_007:sink_channel
	wire          id_router_007_src_ready;                                                                             // rsp_xbar_demux_007:sink_ready -> id_router_007:src_ready
	wire          cmd_xbar_mux_008_src_endofpacket;                                                                    // cmd_xbar_mux_008:src_endofpacket -> burst_adapter_006:sink0_endofpacket
	wire          cmd_xbar_mux_008_src_valid;                                                                          // cmd_xbar_mux_008:src_valid -> burst_adapter_006:sink0_valid
	wire          cmd_xbar_mux_008_src_startofpacket;                                                                  // cmd_xbar_mux_008:src_startofpacket -> burst_adapter_006:sink0_startofpacket
	wire  [112:0] cmd_xbar_mux_008_src_data;                                                                           // cmd_xbar_mux_008:src_data -> burst_adapter_006:sink0_data
	wire    [7:0] cmd_xbar_mux_008_src_channel;                                                                        // cmd_xbar_mux_008:src_channel -> burst_adapter_006:sink0_channel
	wire          cmd_xbar_mux_008_src_ready;                                                                          // burst_adapter_006:sink0_ready -> cmd_xbar_mux_008:src_ready
	wire          id_router_008_src_endofpacket;                                                                       // id_router_008:src_endofpacket -> rsp_xbar_demux_008:sink_endofpacket
	wire          id_router_008_src_valid;                                                                             // id_router_008:src_valid -> rsp_xbar_demux_008:sink_valid
	wire          id_router_008_src_startofpacket;                                                                     // id_router_008:src_startofpacket -> rsp_xbar_demux_008:sink_startofpacket
	wire  [112:0] id_router_008_src_data;                                                                              // id_router_008:src_data -> rsp_xbar_demux_008:sink_data
	wire    [7:0] id_router_008_src_channel;                                                                           // id_router_008:src_channel -> rsp_xbar_demux_008:sink_channel
	wire          id_router_008_src_ready;                                                                             // rsp_xbar_demux_008:sink_ready -> id_router_008:src_ready
	wire          cmd_xbar_mux_009_src_endofpacket;                                                                    // cmd_xbar_mux_009:src_endofpacket -> burst_adapter_007:sink0_endofpacket
	wire          cmd_xbar_mux_009_src_valid;                                                                          // cmd_xbar_mux_009:src_valid -> burst_adapter_007:sink0_valid
	wire          cmd_xbar_mux_009_src_startofpacket;                                                                  // cmd_xbar_mux_009:src_startofpacket -> burst_adapter_007:sink0_startofpacket
	wire  [112:0] cmd_xbar_mux_009_src_data;                                                                           // cmd_xbar_mux_009:src_data -> burst_adapter_007:sink0_data
	wire    [7:0] cmd_xbar_mux_009_src_channel;                                                                        // cmd_xbar_mux_009:src_channel -> burst_adapter_007:sink0_channel
	wire          cmd_xbar_mux_009_src_ready;                                                                          // burst_adapter_007:sink0_ready -> cmd_xbar_mux_009:src_ready
	wire          id_router_009_src_endofpacket;                                                                       // id_router_009:src_endofpacket -> rsp_xbar_demux_009:sink_endofpacket
	wire          id_router_009_src_valid;                                                                             // id_router_009:src_valid -> rsp_xbar_demux_009:sink_valid
	wire          id_router_009_src_startofpacket;                                                                     // id_router_009:src_startofpacket -> rsp_xbar_demux_009:sink_startofpacket
	wire  [112:0] id_router_009_src_data;                                                                              // id_router_009:src_data -> rsp_xbar_demux_009:sink_data
	wire    [7:0] id_router_009_src_channel;                                                                           // id_router_009:src_channel -> rsp_xbar_demux_009:sink_channel
	wire          id_router_009_src_ready;                                                                             // rsp_xbar_demux_009:sink_ready -> id_router_009:src_ready
	wire          cmd_xbar_demux_003_src0_endofpacket;                                                                 // cmd_xbar_demux_003:src0_endofpacket -> cmd_xbar_mux_010:sink0_endofpacket
	wire          cmd_xbar_demux_003_src0_valid;                                                                       // cmd_xbar_demux_003:src0_valid -> cmd_xbar_mux_010:sink0_valid
	wire          cmd_xbar_demux_003_src0_startofpacket;                                                               // cmd_xbar_demux_003:src0_startofpacket -> cmd_xbar_mux_010:sink0_startofpacket
	wire  [233:0] cmd_xbar_demux_003_src0_data;                                                                        // cmd_xbar_demux_003:src0_data -> cmd_xbar_mux_010:sink0_data
	wire    [2:0] cmd_xbar_demux_003_src0_channel;                                                                     // cmd_xbar_demux_003:src0_channel -> cmd_xbar_mux_010:sink0_channel
	wire          cmd_xbar_demux_003_src0_ready;                                                                       // cmd_xbar_mux_010:sink0_ready -> cmd_xbar_demux_003:src0_ready
	wire          cmd_xbar_demux_004_src0_endofpacket;                                                                 // cmd_xbar_demux_004:src0_endofpacket -> cmd_xbar_mux_010:sink1_endofpacket
	wire          cmd_xbar_demux_004_src0_valid;                                                                       // cmd_xbar_demux_004:src0_valid -> cmd_xbar_mux_010:sink1_valid
	wire          cmd_xbar_demux_004_src0_startofpacket;                                                               // cmd_xbar_demux_004:src0_startofpacket -> cmd_xbar_mux_010:sink1_startofpacket
	wire  [233:0] cmd_xbar_demux_004_src0_data;                                                                        // cmd_xbar_demux_004:src0_data -> cmd_xbar_mux_010:sink1_data
	wire    [2:0] cmd_xbar_demux_004_src0_channel;                                                                     // cmd_xbar_demux_004:src0_channel -> cmd_xbar_mux_010:sink1_channel
	wire          cmd_xbar_demux_004_src0_ready;                                                                       // cmd_xbar_mux_010:sink1_ready -> cmd_xbar_demux_004:src0_ready
	wire          cmd_xbar_demux_005_src0_endofpacket;                                                                 // cmd_xbar_demux_005:src0_endofpacket -> cmd_xbar_mux_010:sink2_endofpacket
	wire          cmd_xbar_demux_005_src0_valid;                                                                       // cmd_xbar_demux_005:src0_valid -> cmd_xbar_mux_010:sink2_valid
	wire          cmd_xbar_demux_005_src0_startofpacket;                                                               // cmd_xbar_demux_005:src0_startofpacket -> cmd_xbar_mux_010:sink2_startofpacket
	wire  [233:0] cmd_xbar_demux_005_src0_data;                                                                        // cmd_xbar_demux_005:src0_data -> cmd_xbar_mux_010:sink2_data
	wire    [2:0] cmd_xbar_demux_005_src0_channel;                                                                     // cmd_xbar_demux_005:src0_channel -> cmd_xbar_mux_010:sink2_channel
	wire          cmd_xbar_demux_005_src0_ready;                                                                       // cmd_xbar_mux_010:sink2_ready -> cmd_xbar_demux_005:src0_ready
	wire          rsp_xbar_demux_010_src0_endofpacket;                                                                 // rsp_xbar_demux_010:src0_endofpacket -> hps_0_h2f_axi_master_agent:write_rp_endofpacket
	wire          rsp_xbar_demux_010_src0_valid;                                                                       // rsp_xbar_demux_010:src0_valid -> hps_0_h2f_axi_master_agent:write_rp_valid
	wire          rsp_xbar_demux_010_src0_startofpacket;                                                               // rsp_xbar_demux_010:src0_startofpacket -> hps_0_h2f_axi_master_agent:write_rp_startofpacket
	wire  [233:0] rsp_xbar_demux_010_src0_data;                                                                        // rsp_xbar_demux_010:src0_data -> hps_0_h2f_axi_master_agent:write_rp_data
	wire    [2:0] rsp_xbar_demux_010_src0_channel;                                                                     // rsp_xbar_demux_010:src0_channel -> hps_0_h2f_axi_master_agent:write_rp_channel
	wire          rsp_xbar_demux_010_src1_endofpacket;                                                                 // rsp_xbar_demux_010:src1_endofpacket -> hps_0_h2f_axi_master_agent:read_rp_endofpacket
	wire          rsp_xbar_demux_010_src1_valid;                                                                       // rsp_xbar_demux_010:src1_valid -> hps_0_h2f_axi_master_agent:read_rp_valid
	wire          rsp_xbar_demux_010_src1_startofpacket;                                                               // rsp_xbar_demux_010:src1_startofpacket -> hps_0_h2f_axi_master_agent:read_rp_startofpacket
	wire  [233:0] rsp_xbar_demux_010_src1_data;                                                                        // rsp_xbar_demux_010:src1_data -> hps_0_h2f_axi_master_agent:read_rp_data
	wire    [2:0] rsp_xbar_demux_010_src1_channel;                                                                     // rsp_xbar_demux_010:src1_channel -> hps_0_h2f_axi_master_agent:read_rp_channel
	wire          rsp_xbar_demux_010_src2_endofpacket;                                                                 // rsp_xbar_demux_010:src2_endofpacket -> width_adapter_002:rsp_in_endofpacket
	wire          rsp_xbar_demux_010_src2_valid;                                                                       // rsp_xbar_demux_010:src2_valid -> width_adapter_002:rsp_in_valid
	wire          rsp_xbar_demux_010_src2_startofpacket;                                                               // rsp_xbar_demux_010:src2_startofpacket -> width_adapter_002:rsp_in_startofpacket
	wire  [233:0] rsp_xbar_demux_010_src2_data;                                                                        // rsp_xbar_demux_010:src2_data -> width_adapter_002:rsp_in_data
	wire    [2:0] rsp_xbar_demux_010_src2_channel;                                                                     // rsp_xbar_demux_010:src2_channel -> width_adapter_002:rsp_in_channel
	wire          addr_router_003_src_endofpacket;                                                                     // addr_router_003:src_endofpacket -> cmd_xbar_demux_003:sink_endofpacket
	wire          addr_router_003_src_valid;                                                                           // addr_router_003:src_valid -> cmd_xbar_demux_003:sink_valid
	wire          addr_router_003_src_startofpacket;                                                                   // addr_router_003:src_startofpacket -> cmd_xbar_demux_003:sink_startofpacket
	wire  [233:0] addr_router_003_src_data;                                                                            // addr_router_003:src_data -> cmd_xbar_demux_003:sink_data
	wire    [2:0] addr_router_003_src_channel;                                                                         // addr_router_003:src_channel -> cmd_xbar_demux_003:sink_channel
	wire          addr_router_003_src_ready;                                                                           // cmd_xbar_demux_003:sink_ready -> addr_router_003:src_ready
	wire          rsp_xbar_demux_010_src0_ready;                                                                       // hps_0_h2f_axi_master_agent:write_rp_ready -> rsp_xbar_demux_010:src0_ready
	wire          addr_router_004_src_endofpacket;                                                                     // addr_router_004:src_endofpacket -> cmd_xbar_demux_004:sink_endofpacket
	wire          addr_router_004_src_valid;                                                                           // addr_router_004:src_valid -> cmd_xbar_demux_004:sink_valid
	wire          addr_router_004_src_startofpacket;                                                                   // addr_router_004:src_startofpacket -> cmd_xbar_demux_004:sink_startofpacket
	wire  [233:0] addr_router_004_src_data;                                                                            // addr_router_004:src_data -> cmd_xbar_demux_004:sink_data
	wire    [2:0] addr_router_004_src_channel;                                                                         // addr_router_004:src_channel -> cmd_xbar_demux_004:sink_channel
	wire          addr_router_004_src_ready;                                                                           // cmd_xbar_demux_004:sink_ready -> addr_router_004:src_ready
	wire          rsp_xbar_demux_010_src1_ready;                                                                       // hps_0_h2f_axi_master_agent:read_rp_ready -> rsp_xbar_demux_010:src1_ready
	wire          width_adapter_002_cmd_source_endofpacket;                                                            // width_adapter_002:cmd_out_endofpacket -> cmd_xbar_demux_005:sink_endofpacket
	wire          width_adapter_002_cmd_source_valid;                                                                  // width_adapter_002:cmd_out_valid -> cmd_xbar_demux_005:sink_valid
	wire          width_adapter_002_cmd_source_startofpacket;                                                          // width_adapter_002:cmd_out_startofpacket -> cmd_xbar_demux_005:sink_startofpacket
	wire  [233:0] width_adapter_002_cmd_source_data;                                                                   // width_adapter_002:cmd_out_data -> cmd_xbar_demux_005:sink_data
	wire    [2:0] width_adapter_002_cmd_source_channel;                                                                // width_adapter_002:cmd_out_channel -> cmd_xbar_demux_005:sink_channel
	wire          width_adapter_002_cmd_source_ready;                                                                  // cmd_xbar_demux_005:sink_ready -> width_adapter_002:cmd_out_ready
	wire          rsp_xbar_demux_010_src2_ready;                                                                       // width_adapter_002:rsp_in_ready -> rsp_xbar_demux_010:src2_ready
	wire          cmd_xbar_mux_010_src_endofpacket;                                                                    // cmd_xbar_mux_010:src_endofpacket -> width_adapter_003:cmd_in_endofpacket
	wire          cmd_xbar_mux_010_src_valid;                                                                          // cmd_xbar_mux_010:src_valid -> width_adapter_003:cmd_in_valid
	wire          cmd_xbar_mux_010_src_startofpacket;                                                                  // cmd_xbar_mux_010:src_startofpacket -> width_adapter_003:cmd_in_startofpacket
	wire  [233:0] cmd_xbar_mux_010_src_data;                                                                           // cmd_xbar_mux_010:src_data -> width_adapter_003:cmd_in_data
	wire    [2:0] cmd_xbar_mux_010_src_channel;                                                                        // cmd_xbar_mux_010:src_channel -> width_adapter_003:cmd_in_channel
	wire          cmd_xbar_mux_010_src_ready;                                                                          // width_adapter_003:cmd_in_ready -> cmd_xbar_mux_010:src_ready
	wire          width_adapter_003_rsp_source_endofpacket;                                                            // width_adapter_003:rsp_out_endofpacket -> rsp_xbar_demux_010:sink_endofpacket
	wire          width_adapter_003_rsp_source_valid;                                                                  // width_adapter_003:rsp_out_valid -> rsp_xbar_demux_010:sink_valid
	wire          width_adapter_003_rsp_source_startofpacket;                                                          // width_adapter_003:rsp_out_startofpacket -> rsp_xbar_demux_010:sink_startofpacket
	wire  [233:0] width_adapter_003_rsp_source_data;                                                                   // width_adapter_003:rsp_out_data -> rsp_xbar_demux_010:sink_data
	wire    [2:0] width_adapter_003_rsp_source_channel;                                                                // width_adapter_003:rsp_out_channel -> rsp_xbar_demux_010:sink_channel
	wire          width_adapter_003_rsp_source_ready;                                                                  // rsp_xbar_demux_010:sink_ready -> width_adapter_003:rsp_out_ready
	wire          crosser_out_endofpacket;                                                                             // crosser:out_endofpacket -> cmd_xbar_mux_007:sink0_endofpacket
	wire          crosser_out_valid;                                                                                   // crosser:out_valid -> cmd_xbar_mux_007:sink0_valid
	wire          crosser_out_startofpacket;                                                                           // crosser:out_startofpacket -> cmd_xbar_mux_007:sink0_startofpacket
	wire  [112:0] crosser_out_data;                                                                                    // crosser:out_data -> cmd_xbar_mux_007:sink0_data
	wire    [7:0] crosser_out_channel;                                                                                 // crosser:out_channel -> cmd_xbar_mux_007:sink0_channel
	wire          crosser_out_ready;                                                                                   // cmd_xbar_mux_007:sink0_ready -> crosser:out_ready
	wire          cmd_xbar_demux_001_src5_endofpacket;                                                                 // cmd_xbar_demux_001:src5_endofpacket -> crosser:in_endofpacket
	wire          cmd_xbar_demux_001_src5_valid;                                                                       // cmd_xbar_demux_001:src5_valid -> crosser:in_valid
	wire          cmd_xbar_demux_001_src5_startofpacket;                                                               // cmd_xbar_demux_001:src5_startofpacket -> crosser:in_startofpacket
	wire  [112:0] cmd_xbar_demux_001_src5_data;                                                                        // cmd_xbar_demux_001:src5_data -> crosser:in_data
	wire    [7:0] cmd_xbar_demux_001_src5_channel;                                                                     // cmd_xbar_demux_001:src5_channel -> crosser:in_channel
	wire          cmd_xbar_demux_001_src5_ready;                                                                       // crosser:in_ready -> cmd_xbar_demux_001:src5_ready
	wire          crosser_001_out_endofpacket;                                                                         // crosser_001:out_endofpacket -> cmd_xbar_mux_008:sink0_endofpacket
	wire          crosser_001_out_valid;                                                                               // crosser_001:out_valid -> cmd_xbar_mux_008:sink0_valid
	wire          crosser_001_out_startofpacket;                                                                       // crosser_001:out_startofpacket -> cmd_xbar_mux_008:sink0_startofpacket
	wire  [112:0] crosser_001_out_data;                                                                                // crosser_001:out_data -> cmd_xbar_mux_008:sink0_data
	wire    [7:0] crosser_001_out_channel;                                                                             // crosser_001:out_channel -> cmd_xbar_mux_008:sink0_channel
	wire          crosser_001_out_ready;                                                                               // cmd_xbar_mux_008:sink0_ready -> crosser_001:out_ready
	wire          cmd_xbar_demux_001_src6_endofpacket;                                                                 // cmd_xbar_demux_001:src6_endofpacket -> crosser_001:in_endofpacket
	wire          cmd_xbar_demux_001_src6_valid;                                                                       // cmd_xbar_demux_001:src6_valid -> crosser_001:in_valid
	wire          cmd_xbar_demux_001_src6_startofpacket;                                                               // cmd_xbar_demux_001:src6_startofpacket -> crosser_001:in_startofpacket
	wire  [112:0] cmd_xbar_demux_001_src6_data;                                                                        // cmd_xbar_demux_001:src6_data -> crosser_001:in_data
	wire    [7:0] cmd_xbar_demux_001_src6_channel;                                                                     // cmd_xbar_demux_001:src6_channel -> crosser_001:in_channel
	wire          cmd_xbar_demux_001_src6_ready;                                                                       // crosser_001:in_ready -> cmd_xbar_demux_001:src6_ready
	wire          crosser_002_out_endofpacket;                                                                         // crosser_002:out_endofpacket -> cmd_xbar_mux_009:sink0_endofpacket
	wire          crosser_002_out_valid;                                                                               // crosser_002:out_valid -> cmd_xbar_mux_009:sink0_valid
	wire          crosser_002_out_startofpacket;                                                                       // crosser_002:out_startofpacket -> cmd_xbar_mux_009:sink0_startofpacket
	wire  [112:0] crosser_002_out_data;                                                                                // crosser_002:out_data -> cmd_xbar_mux_009:sink0_data
	wire    [7:0] crosser_002_out_channel;                                                                             // crosser_002:out_channel -> cmd_xbar_mux_009:sink0_channel
	wire          crosser_002_out_ready;                                                                               // cmd_xbar_mux_009:sink0_ready -> crosser_002:out_ready
	wire          cmd_xbar_demux_001_src7_endofpacket;                                                                 // cmd_xbar_demux_001:src7_endofpacket -> crosser_002:in_endofpacket
	wire          cmd_xbar_demux_001_src7_valid;                                                                       // cmd_xbar_demux_001:src7_valid -> crosser_002:in_valid
	wire          cmd_xbar_demux_001_src7_startofpacket;                                                               // cmd_xbar_demux_001:src7_startofpacket -> crosser_002:in_startofpacket
	wire  [112:0] cmd_xbar_demux_001_src7_data;                                                                        // cmd_xbar_demux_001:src7_data -> crosser_002:in_data
	wire    [7:0] cmd_xbar_demux_001_src7_channel;                                                                     // cmd_xbar_demux_001:src7_channel -> crosser_002:in_channel
	wire          cmd_xbar_demux_001_src7_ready;                                                                       // crosser_002:in_ready -> cmd_xbar_demux_001:src7_ready
	wire          crosser_003_out_endofpacket;                                                                         // crosser_003:out_endofpacket -> cmd_xbar_mux_007:sink1_endofpacket
	wire          crosser_003_out_valid;                                                                               // crosser_003:out_valid -> cmd_xbar_mux_007:sink1_valid
	wire          crosser_003_out_startofpacket;                                                                       // crosser_003:out_startofpacket -> cmd_xbar_mux_007:sink1_startofpacket
	wire  [112:0] crosser_003_out_data;                                                                                // crosser_003:out_data -> cmd_xbar_mux_007:sink1_data
	wire    [7:0] crosser_003_out_channel;                                                                             // crosser_003:out_channel -> cmd_xbar_mux_007:sink1_channel
	wire          crosser_003_out_ready;                                                                               // cmd_xbar_mux_007:sink1_ready -> crosser_003:out_ready
	wire          cmd_xbar_demux_002_src5_endofpacket;                                                                 // cmd_xbar_demux_002:src5_endofpacket -> crosser_003:in_endofpacket
	wire          cmd_xbar_demux_002_src5_valid;                                                                       // cmd_xbar_demux_002:src5_valid -> crosser_003:in_valid
	wire          cmd_xbar_demux_002_src5_startofpacket;                                                               // cmd_xbar_demux_002:src5_startofpacket -> crosser_003:in_startofpacket
	wire  [112:0] cmd_xbar_demux_002_src5_data;                                                                        // cmd_xbar_demux_002:src5_data -> crosser_003:in_data
	wire    [7:0] cmd_xbar_demux_002_src5_channel;                                                                     // cmd_xbar_demux_002:src5_channel -> crosser_003:in_channel
	wire          cmd_xbar_demux_002_src5_ready;                                                                       // crosser_003:in_ready -> cmd_xbar_demux_002:src5_ready
	wire          crosser_004_out_endofpacket;                                                                         // crosser_004:out_endofpacket -> cmd_xbar_mux_008:sink1_endofpacket
	wire          crosser_004_out_valid;                                                                               // crosser_004:out_valid -> cmd_xbar_mux_008:sink1_valid
	wire          crosser_004_out_startofpacket;                                                                       // crosser_004:out_startofpacket -> cmd_xbar_mux_008:sink1_startofpacket
	wire  [112:0] crosser_004_out_data;                                                                                // crosser_004:out_data -> cmd_xbar_mux_008:sink1_data
	wire    [7:0] crosser_004_out_channel;                                                                             // crosser_004:out_channel -> cmd_xbar_mux_008:sink1_channel
	wire          crosser_004_out_ready;                                                                               // cmd_xbar_mux_008:sink1_ready -> crosser_004:out_ready
	wire          cmd_xbar_demux_002_src6_endofpacket;                                                                 // cmd_xbar_demux_002:src6_endofpacket -> crosser_004:in_endofpacket
	wire          cmd_xbar_demux_002_src6_valid;                                                                       // cmd_xbar_demux_002:src6_valid -> crosser_004:in_valid
	wire          cmd_xbar_demux_002_src6_startofpacket;                                                               // cmd_xbar_demux_002:src6_startofpacket -> crosser_004:in_startofpacket
	wire  [112:0] cmd_xbar_demux_002_src6_data;                                                                        // cmd_xbar_demux_002:src6_data -> crosser_004:in_data
	wire    [7:0] cmd_xbar_demux_002_src6_channel;                                                                     // cmd_xbar_demux_002:src6_channel -> crosser_004:in_channel
	wire          cmd_xbar_demux_002_src6_ready;                                                                       // crosser_004:in_ready -> cmd_xbar_demux_002:src6_ready
	wire          crosser_005_out_endofpacket;                                                                         // crosser_005:out_endofpacket -> cmd_xbar_mux_009:sink1_endofpacket
	wire          crosser_005_out_valid;                                                                               // crosser_005:out_valid -> cmd_xbar_mux_009:sink1_valid
	wire          crosser_005_out_startofpacket;                                                                       // crosser_005:out_startofpacket -> cmd_xbar_mux_009:sink1_startofpacket
	wire  [112:0] crosser_005_out_data;                                                                                // crosser_005:out_data -> cmd_xbar_mux_009:sink1_data
	wire    [7:0] crosser_005_out_channel;                                                                             // crosser_005:out_channel -> cmd_xbar_mux_009:sink1_channel
	wire          crosser_005_out_ready;                                                                               // cmd_xbar_mux_009:sink1_ready -> crosser_005:out_ready
	wire          cmd_xbar_demux_002_src7_endofpacket;                                                                 // cmd_xbar_demux_002:src7_endofpacket -> crosser_005:in_endofpacket
	wire          cmd_xbar_demux_002_src7_valid;                                                                       // cmd_xbar_demux_002:src7_valid -> crosser_005:in_valid
	wire          cmd_xbar_demux_002_src7_startofpacket;                                                               // cmd_xbar_demux_002:src7_startofpacket -> crosser_005:in_startofpacket
	wire  [112:0] cmd_xbar_demux_002_src7_data;                                                                        // cmd_xbar_demux_002:src7_data -> crosser_005:in_data
	wire    [7:0] cmd_xbar_demux_002_src7_channel;                                                                     // cmd_xbar_demux_002:src7_channel -> crosser_005:in_channel
	wire          cmd_xbar_demux_002_src7_ready;                                                                       // crosser_005:in_ready -> cmd_xbar_demux_002:src7_ready
	wire          crosser_006_out_endofpacket;                                                                         // crosser_006:out_endofpacket -> rsp_xbar_mux_001:sink5_endofpacket
	wire          crosser_006_out_valid;                                                                               // crosser_006:out_valid -> rsp_xbar_mux_001:sink5_valid
	wire          crosser_006_out_startofpacket;                                                                       // crosser_006:out_startofpacket -> rsp_xbar_mux_001:sink5_startofpacket
	wire  [112:0] crosser_006_out_data;                                                                                // crosser_006:out_data -> rsp_xbar_mux_001:sink5_data
	wire    [7:0] crosser_006_out_channel;                                                                             // crosser_006:out_channel -> rsp_xbar_mux_001:sink5_channel
	wire          crosser_006_out_ready;                                                                               // rsp_xbar_mux_001:sink5_ready -> crosser_006:out_ready
	wire          rsp_xbar_demux_007_src0_endofpacket;                                                                 // rsp_xbar_demux_007:src0_endofpacket -> crosser_006:in_endofpacket
	wire          rsp_xbar_demux_007_src0_valid;                                                                       // rsp_xbar_demux_007:src0_valid -> crosser_006:in_valid
	wire          rsp_xbar_demux_007_src0_startofpacket;                                                               // rsp_xbar_demux_007:src0_startofpacket -> crosser_006:in_startofpacket
	wire  [112:0] rsp_xbar_demux_007_src0_data;                                                                        // rsp_xbar_demux_007:src0_data -> crosser_006:in_data
	wire    [7:0] rsp_xbar_demux_007_src0_channel;                                                                     // rsp_xbar_demux_007:src0_channel -> crosser_006:in_channel
	wire          rsp_xbar_demux_007_src0_ready;                                                                       // crosser_006:in_ready -> rsp_xbar_demux_007:src0_ready
	wire          crosser_007_out_endofpacket;                                                                         // crosser_007:out_endofpacket -> rsp_xbar_mux_002:sink5_endofpacket
	wire          crosser_007_out_valid;                                                                               // crosser_007:out_valid -> rsp_xbar_mux_002:sink5_valid
	wire          crosser_007_out_startofpacket;                                                                       // crosser_007:out_startofpacket -> rsp_xbar_mux_002:sink5_startofpacket
	wire  [112:0] crosser_007_out_data;                                                                                // crosser_007:out_data -> rsp_xbar_mux_002:sink5_data
	wire    [7:0] crosser_007_out_channel;                                                                             // crosser_007:out_channel -> rsp_xbar_mux_002:sink5_channel
	wire          crosser_007_out_ready;                                                                               // rsp_xbar_mux_002:sink5_ready -> crosser_007:out_ready
	wire          rsp_xbar_demux_007_src1_endofpacket;                                                                 // rsp_xbar_demux_007:src1_endofpacket -> crosser_007:in_endofpacket
	wire          rsp_xbar_demux_007_src1_valid;                                                                       // rsp_xbar_demux_007:src1_valid -> crosser_007:in_valid
	wire          rsp_xbar_demux_007_src1_startofpacket;                                                               // rsp_xbar_demux_007:src1_startofpacket -> crosser_007:in_startofpacket
	wire  [112:0] rsp_xbar_demux_007_src1_data;                                                                        // rsp_xbar_demux_007:src1_data -> crosser_007:in_data
	wire    [7:0] rsp_xbar_demux_007_src1_channel;                                                                     // rsp_xbar_demux_007:src1_channel -> crosser_007:in_channel
	wire          rsp_xbar_demux_007_src1_ready;                                                                       // crosser_007:in_ready -> rsp_xbar_demux_007:src1_ready
	wire          crosser_008_out_endofpacket;                                                                         // crosser_008:out_endofpacket -> rsp_xbar_mux_001:sink6_endofpacket
	wire          crosser_008_out_valid;                                                                               // crosser_008:out_valid -> rsp_xbar_mux_001:sink6_valid
	wire          crosser_008_out_startofpacket;                                                                       // crosser_008:out_startofpacket -> rsp_xbar_mux_001:sink6_startofpacket
	wire  [112:0] crosser_008_out_data;                                                                                // crosser_008:out_data -> rsp_xbar_mux_001:sink6_data
	wire    [7:0] crosser_008_out_channel;                                                                             // crosser_008:out_channel -> rsp_xbar_mux_001:sink6_channel
	wire          crosser_008_out_ready;                                                                               // rsp_xbar_mux_001:sink6_ready -> crosser_008:out_ready
	wire          rsp_xbar_demux_008_src0_endofpacket;                                                                 // rsp_xbar_demux_008:src0_endofpacket -> crosser_008:in_endofpacket
	wire          rsp_xbar_demux_008_src0_valid;                                                                       // rsp_xbar_demux_008:src0_valid -> crosser_008:in_valid
	wire          rsp_xbar_demux_008_src0_startofpacket;                                                               // rsp_xbar_demux_008:src0_startofpacket -> crosser_008:in_startofpacket
	wire  [112:0] rsp_xbar_demux_008_src0_data;                                                                        // rsp_xbar_demux_008:src0_data -> crosser_008:in_data
	wire    [7:0] rsp_xbar_demux_008_src0_channel;                                                                     // rsp_xbar_demux_008:src0_channel -> crosser_008:in_channel
	wire          rsp_xbar_demux_008_src0_ready;                                                                       // crosser_008:in_ready -> rsp_xbar_demux_008:src0_ready
	wire          crosser_009_out_endofpacket;                                                                         // crosser_009:out_endofpacket -> rsp_xbar_mux_002:sink6_endofpacket
	wire          crosser_009_out_valid;                                                                               // crosser_009:out_valid -> rsp_xbar_mux_002:sink6_valid
	wire          crosser_009_out_startofpacket;                                                                       // crosser_009:out_startofpacket -> rsp_xbar_mux_002:sink6_startofpacket
	wire  [112:0] crosser_009_out_data;                                                                                // crosser_009:out_data -> rsp_xbar_mux_002:sink6_data
	wire    [7:0] crosser_009_out_channel;                                                                             // crosser_009:out_channel -> rsp_xbar_mux_002:sink6_channel
	wire          crosser_009_out_ready;                                                                               // rsp_xbar_mux_002:sink6_ready -> crosser_009:out_ready
	wire          rsp_xbar_demux_008_src1_endofpacket;                                                                 // rsp_xbar_demux_008:src1_endofpacket -> crosser_009:in_endofpacket
	wire          rsp_xbar_demux_008_src1_valid;                                                                       // rsp_xbar_demux_008:src1_valid -> crosser_009:in_valid
	wire          rsp_xbar_demux_008_src1_startofpacket;                                                               // rsp_xbar_demux_008:src1_startofpacket -> crosser_009:in_startofpacket
	wire  [112:0] rsp_xbar_demux_008_src1_data;                                                                        // rsp_xbar_demux_008:src1_data -> crosser_009:in_data
	wire    [7:0] rsp_xbar_demux_008_src1_channel;                                                                     // rsp_xbar_demux_008:src1_channel -> crosser_009:in_channel
	wire          rsp_xbar_demux_008_src1_ready;                                                                       // crosser_009:in_ready -> rsp_xbar_demux_008:src1_ready
	wire          crosser_010_out_endofpacket;                                                                         // crosser_010:out_endofpacket -> rsp_xbar_mux_001:sink7_endofpacket
	wire          crosser_010_out_valid;                                                                               // crosser_010:out_valid -> rsp_xbar_mux_001:sink7_valid
	wire          crosser_010_out_startofpacket;                                                                       // crosser_010:out_startofpacket -> rsp_xbar_mux_001:sink7_startofpacket
	wire  [112:0] crosser_010_out_data;                                                                                // crosser_010:out_data -> rsp_xbar_mux_001:sink7_data
	wire    [7:0] crosser_010_out_channel;                                                                             // crosser_010:out_channel -> rsp_xbar_mux_001:sink7_channel
	wire          crosser_010_out_ready;                                                                               // rsp_xbar_mux_001:sink7_ready -> crosser_010:out_ready
	wire          rsp_xbar_demux_009_src0_endofpacket;                                                                 // rsp_xbar_demux_009:src0_endofpacket -> crosser_010:in_endofpacket
	wire          rsp_xbar_demux_009_src0_valid;                                                                       // rsp_xbar_demux_009:src0_valid -> crosser_010:in_valid
	wire          rsp_xbar_demux_009_src0_startofpacket;                                                               // rsp_xbar_demux_009:src0_startofpacket -> crosser_010:in_startofpacket
	wire  [112:0] rsp_xbar_demux_009_src0_data;                                                                        // rsp_xbar_demux_009:src0_data -> crosser_010:in_data
	wire    [7:0] rsp_xbar_demux_009_src0_channel;                                                                     // rsp_xbar_demux_009:src0_channel -> crosser_010:in_channel
	wire          rsp_xbar_demux_009_src0_ready;                                                                       // crosser_010:in_ready -> rsp_xbar_demux_009:src0_ready
	wire          crosser_011_out_endofpacket;                                                                         // crosser_011:out_endofpacket -> rsp_xbar_mux_002:sink7_endofpacket
	wire          crosser_011_out_valid;                                                                               // crosser_011:out_valid -> rsp_xbar_mux_002:sink7_valid
	wire          crosser_011_out_startofpacket;                                                                       // crosser_011:out_startofpacket -> rsp_xbar_mux_002:sink7_startofpacket
	wire  [112:0] crosser_011_out_data;                                                                                // crosser_011:out_data -> rsp_xbar_mux_002:sink7_data
	wire    [7:0] crosser_011_out_channel;                                                                             // crosser_011:out_channel -> rsp_xbar_mux_002:sink7_channel
	wire          crosser_011_out_ready;                                                                               // rsp_xbar_mux_002:sink7_ready -> crosser_011:out_ready
	wire          rsp_xbar_demux_009_src1_endofpacket;                                                                 // rsp_xbar_demux_009:src1_endofpacket -> crosser_011:in_endofpacket
	wire          rsp_xbar_demux_009_src1_valid;                                                                       // rsp_xbar_demux_009:src1_valid -> crosser_011:in_valid
	wire          rsp_xbar_demux_009_src1_startofpacket;                                                               // rsp_xbar_demux_009:src1_startofpacket -> crosser_011:in_startofpacket
	wire  [112:0] rsp_xbar_demux_009_src1_data;                                                                        // rsp_xbar_demux_009:src1_data -> crosser_011:in_data
	wire    [7:0] rsp_xbar_demux_009_src1_channel;                                                                     // rsp_xbar_demux_009:src1_channel -> crosser_011:in_channel
	wire          rsp_xbar_demux_009_src1_ready;                                                                       // crosser_011:in_ready -> rsp_xbar_demux_009:src1_ready
	wire    [1:0] limiter_cmd_valid_data;                                                                              // limiter:cmd_src_valid -> cmd_xbar_demux:sink_valid
	wire    [7:0] limiter_001_cmd_valid_data;                                                                          // limiter_001:cmd_src_valid -> cmd_xbar_demux_001:sink_valid
	wire    [7:0] limiter_002_cmd_valid_data;                                                                          // limiter_002:cmd_src_valid -> cmd_xbar_demux_002:sink_valid
	wire          irq_mapper_receiver0_irq;                                                                            // jtag_uart:av_irq -> irq_mapper:receiver0_irq
	wire          irq_mapper_receiver1_irq;                                                                            // button_pio:irq -> irq_mapper:receiver1_irq
	wire          irq_mapper_receiver2_irq;                                                                            // dipsw_pio:irq -> irq_mapper:receiver2_irq
	wire   [31:0] hps_0_f2h_irq0_irq;                                                                                  // irq_mapper:sender_irq -> hps_0:f2h_irq_p0
	wire   [31:0] hps_0_f2h_irq1_irq;                                                                                  // irq_mapper_001:sender_irq -> hps_0:f2h_irq_p1
	wire          log_generate_0_dout_endofpacket;                                                                     // LOG_Generate_0:dout_eop -> avalon_st_adapter:in_0_endofpacket
	wire          log_generate_0_dout_valid;                                                                           // LOG_Generate_0:dout_valid -> avalon_st_adapter:in_0_valid
	wire          log_generate_0_dout_startofpacket;                                                                   // LOG_Generate_0:dout_sop -> avalon_st_adapter:in_0_startofpacket
	wire    [1:0] log_generate_0_dout_empty;                                                                           // LOG_Generate_0:dout_empty -> avalon_st_adapter:in_0_empty
	wire   [23:0] log_generate_0_dout_data;                                                                            // LOG_Generate_0:dout_data -> avalon_st_adapter:in_0_data
	wire          log_generate_0_dout_ready;                                                                           // avalon_st_adapter:in_0_ready -> LOG_Generate_0:dout_ready
	wire          avalon_st_adapter_out_0_endofpacket;                                                                 // avalon_st_adapter:out_0_endofpacket -> timing_adapter_0:in_endofpacket
	wire          avalon_st_adapter_out_0_valid;                                                                       // avalon_st_adapter:out_0_valid -> timing_adapter_0:in_valid
	wire          avalon_st_adapter_out_0_startofpacket;                                                               // avalon_st_adapter:out_0_startofpacket -> timing_adapter_0:in_startofpacket
	wire   [23:0] avalon_st_adapter_out_0_data;                                                                        // avalon_st_adapter:out_0_data -> timing_adapter_0:in_data
	wire          avalon_st_adapter_out_0_ready;                                                                       // timing_adapter_0:in_ready -> avalon_st_adapter:out_0_ready

	soc_system_hps_0 #(
		.F2S_Width (2),
		.S2F_Width (3)
	) hps_0 (
		.mem_a                    (memory_mem_a),                                        //            memory.mem_a
		.mem_ba                   (memory_mem_ba),                                       //                  .mem_ba
		.mem_ck                   (memory_mem_ck),                                       //                  .mem_ck
		.mem_ck_n                 (memory_mem_ck_n),                                     //                  .mem_ck_n
		.mem_cke                  (memory_mem_cke),                                      //                  .mem_cke
		.mem_cs_n                 (memory_mem_cs_n),                                     //                  .mem_cs_n
		.mem_ras_n                (memory_mem_ras_n),                                    //                  .mem_ras_n
		.mem_cas_n                (memory_mem_cas_n),                                    //                  .mem_cas_n
		.mem_we_n                 (memory_mem_we_n),                                     //                  .mem_we_n
		.mem_reset_n              (memory_mem_reset_n),                                  //                  .mem_reset_n
		.mem_dq                   (memory_mem_dq),                                       //                  .mem_dq
		.mem_dqs                  (memory_mem_dqs),                                      //                  .mem_dqs
		.mem_dqs_n                (memory_mem_dqs_n),                                    //                  .mem_dqs_n
		.mem_odt                  (memory_mem_odt),                                      //                  .mem_odt
		.mem_dm                   (memory_mem_dm),                                       //                  .mem_dm
		.oct_rzqin                (memory_oct_rzqin),                                    //                  .oct_rzqin
		.hps_io_emac1_inst_TX_CLK (hps_0_hps_io_hps_io_emac1_inst_TX_CLK),               //            hps_io.hps_io_emac1_inst_TX_CLK
		.hps_io_emac1_inst_TXD0   (hps_0_hps_io_hps_io_emac1_inst_TXD0),                 //                  .hps_io_emac1_inst_TXD0
		.hps_io_emac1_inst_TXD1   (hps_0_hps_io_hps_io_emac1_inst_TXD1),                 //                  .hps_io_emac1_inst_TXD1
		.hps_io_emac1_inst_TXD2   (hps_0_hps_io_hps_io_emac1_inst_TXD2),                 //                  .hps_io_emac1_inst_TXD2
		.hps_io_emac1_inst_TXD3   (hps_0_hps_io_hps_io_emac1_inst_TXD3),                 //                  .hps_io_emac1_inst_TXD3
		.hps_io_emac1_inst_RXD0   (hps_0_hps_io_hps_io_emac1_inst_RXD0),                 //                  .hps_io_emac1_inst_RXD0
		.hps_io_emac1_inst_MDIO   (hps_0_hps_io_hps_io_emac1_inst_MDIO),                 //                  .hps_io_emac1_inst_MDIO
		.hps_io_emac1_inst_MDC    (hps_0_hps_io_hps_io_emac1_inst_MDC),                  //                  .hps_io_emac1_inst_MDC
		.hps_io_emac1_inst_RX_CTL (hps_0_hps_io_hps_io_emac1_inst_RX_CTL),               //                  .hps_io_emac1_inst_RX_CTL
		.hps_io_emac1_inst_TX_CTL (hps_0_hps_io_hps_io_emac1_inst_TX_CTL),               //                  .hps_io_emac1_inst_TX_CTL
		.hps_io_emac1_inst_RX_CLK (hps_0_hps_io_hps_io_emac1_inst_RX_CLK),               //                  .hps_io_emac1_inst_RX_CLK
		.hps_io_emac1_inst_RXD1   (hps_0_hps_io_hps_io_emac1_inst_RXD1),                 //                  .hps_io_emac1_inst_RXD1
		.hps_io_emac1_inst_RXD2   (hps_0_hps_io_hps_io_emac1_inst_RXD2),                 //                  .hps_io_emac1_inst_RXD2
		.hps_io_emac1_inst_RXD3   (hps_0_hps_io_hps_io_emac1_inst_RXD3),                 //                  .hps_io_emac1_inst_RXD3
		.hps_io_qspi_inst_IO0     (hps_0_hps_io_hps_io_qspi_inst_IO0),                   //                  .hps_io_qspi_inst_IO0
		.hps_io_qspi_inst_IO1     (hps_0_hps_io_hps_io_qspi_inst_IO1),                   //                  .hps_io_qspi_inst_IO1
		.hps_io_qspi_inst_IO2     (hps_0_hps_io_hps_io_qspi_inst_IO2),                   //                  .hps_io_qspi_inst_IO2
		.hps_io_qspi_inst_IO3     (hps_0_hps_io_hps_io_qspi_inst_IO3),                   //                  .hps_io_qspi_inst_IO3
		.hps_io_qspi_inst_SS0     (hps_0_hps_io_hps_io_qspi_inst_SS0),                   //                  .hps_io_qspi_inst_SS0
		.hps_io_qspi_inst_CLK     (hps_0_hps_io_hps_io_qspi_inst_CLK),                   //                  .hps_io_qspi_inst_CLK
		.hps_io_sdio_inst_CMD     (hps_0_hps_io_hps_io_sdio_inst_CMD),                   //                  .hps_io_sdio_inst_CMD
		.hps_io_sdio_inst_D0      (hps_0_hps_io_hps_io_sdio_inst_D0),                    //                  .hps_io_sdio_inst_D0
		.hps_io_sdio_inst_D1      (hps_0_hps_io_hps_io_sdio_inst_D1),                    //                  .hps_io_sdio_inst_D1
		.hps_io_sdio_inst_CLK     (hps_0_hps_io_hps_io_sdio_inst_CLK),                   //                  .hps_io_sdio_inst_CLK
		.hps_io_sdio_inst_D2      (hps_0_hps_io_hps_io_sdio_inst_D2),                    //                  .hps_io_sdio_inst_D2
		.hps_io_sdio_inst_D3      (hps_0_hps_io_hps_io_sdio_inst_D3),                    //                  .hps_io_sdio_inst_D3
		.hps_io_usb1_inst_D0      (hps_0_hps_io_hps_io_usb1_inst_D0),                    //                  .hps_io_usb1_inst_D0
		.hps_io_usb1_inst_D1      (hps_0_hps_io_hps_io_usb1_inst_D1),                    //                  .hps_io_usb1_inst_D1
		.hps_io_usb1_inst_D2      (hps_0_hps_io_hps_io_usb1_inst_D2),                    //                  .hps_io_usb1_inst_D2
		.hps_io_usb1_inst_D3      (hps_0_hps_io_hps_io_usb1_inst_D3),                    //                  .hps_io_usb1_inst_D3
		.hps_io_usb1_inst_D4      (hps_0_hps_io_hps_io_usb1_inst_D4),                    //                  .hps_io_usb1_inst_D4
		.hps_io_usb1_inst_D5      (hps_0_hps_io_hps_io_usb1_inst_D5),                    //                  .hps_io_usb1_inst_D5
		.hps_io_usb1_inst_D6      (hps_0_hps_io_hps_io_usb1_inst_D6),                    //                  .hps_io_usb1_inst_D6
		.hps_io_usb1_inst_D7      (hps_0_hps_io_hps_io_usb1_inst_D7),                    //                  .hps_io_usb1_inst_D7
		.hps_io_usb1_inst_CLK     (hps_0_hps_io_hps_io_usb1_inst_CLK),                   //                  .hps_io_usb1_inst_CLK
		.hps_io_usb1_inst_STP     (hps_0_hps_io_hps_io_usb1_inst_STP),                   //                  .hps_io_usb1_inst_STP
		.hps_io_usb1_inst_DIR     (hps_0_hps_io_hps_io_usb1_inst_DIR),                   //                  .hps_io_usb1_inst_DIR
		.hps_io_usb1_inst_NXT     (hps_0_hps_io_hps_io_usb1_inst_NXT),                   //                  .hps_io_usb1_inst_NXT
		.hps_io_spim1_inst_CLK    (hps_0_hps_io_hps_io_spim1_inst_CLK),                  //                  .hps_io_spim1_inst_CLK
		.hps_io_spim1_inst_MOSI   (hps_0_hps_io_hps_io_spim1_inst_MOSI),                 //                  .hps_io_spim1_inst_MOSI
		.hps_io_spim1_inst_MISO   (hps_0_hps_io_hps_io_spim1_inst_MISO),                 //                  .hps_io_spim1_inst_MISO
		.hps_io_spim1_inst_SS0    (hps_0_hps_io_hps_io_spim1_inst_SS0),                  //                  .hps_io_spim1_inst_SS0
		.hps_io_uart0_inst_RX     (hps_0_hps_io_hps_io_uart0_inst_RX),                   //                  .hps_io_uart0_inst_RX
		.hps_io_uart0_inst_TX     (hps_0_hps_io_hps_io_uart0_inst_TX),                   //                  .hps_io_uart0_inst_TX
		.hps_io_i2c0_inst_SDA     (hps_0_hps_io_hps_io_i2c0_inst_SDA),                   //                  .hps_io_i2c0_inst_SDA
		.hps_io_i2c0_inst_SCL     (hps_0_hps_io_hps_io_i2c0_inst_SCL),                   //                  .hps_io_i2c0_inst_SCL
		.hps_io_i2c1_inst_SDA     (hps_0_hps_io_hps_io_i2c1_inst_SDA),                   //                  .hps_io_i2c1_inst_SDA
		.hps_io_i2c1_inst_SCL     (hps_0_hps_io_hps_io_i2c1_inst_SCL),                   //                  .hps_io_i2c1_inst_SCL
		.hps_io_gpio_inst_GPIO09  (hps_0_hps_io_hps_io_gpio_inst_GPIO09),                //                  .hps_io_gpio_inst_GPIO09
		.hps_io_gpio_inst_GPIO35  (hps_0_hps_io_hps_io_gpio_inst_GPIO35),                //                  .hps_io_gpio_inst_GPIO35
		.hps_io_gpio_inst_GPIO40  (hps_0_hps_io_hps_io_gpio_inst_GPIO40),                //                  .hps_io_gpio_inst_GPIO40
		.hps_io_gpio_inst_GPIO41  (hps_0_hps_io_hps_io_gpio_inst_GPIO41),                //                  .hps_io_gpio_inst_GPIO41
		.hps_io_gpio_inst_GPIO48  (hps_0_hps_io_hps_io_gpio_inst_GPIO48),                //                  .hps_io_gpio_inst_GPIO48
		.hps_io_gpio_inst_GPIO53  (hps_0_hps_io_hps_io_gpio_inst_GPIO53),                //                  .hps_io_gpio_inst_GPIO53
		.hps_io_gpio_inst_GPIO54  (hps_0_hps_io_hps_io_gpio_inst_GPIO54),                //                  .hps_io_gpio_inst_GPIO54
		.hps_io_gpio_inst_GPIO61  (hps_0_hps_io_hps_io_gpio_inst_GPIO61),                //                  .hps_io_gpio_inst_GPIO61
		.h2f_rst_n                (hps_0_h2f_reset_reset_n),                             //         h2f_reset.reset_n
		.h2f_axi_clk              (pll_sdram_outclk1_clk),                               //     h2f_axi_clock.clk
		.h2f_AWID                 (hps_0_h2f_axi_master_awid),                           //    h2f_axi_master.awid
		.h2f_AWADDR               (hps_0_h2f_axi_master_awaddr),                         //                  .awaddr
		.h2f_AWLEN                (hps_0_h2f_axi_master_awlen),                          //                  .awlen
		.h2f_AWSIZE               (hps_0_h2f_axi_master_awsize),                         //                  .awsize
		.h2f_AWBURST              (hps_0_h2f_axi_master_awburst),                        //                  .awburst
		.h2f_AWLOCK               (hps_0_h2f_axi_master_awlock),                         //                  .awlock
		.h2f_AWCACHE              (hps_0_h2f_axi_master_awcache),                        //                  .awcache
		.h2f_AWPROT               (hps_0_h2f_axi_master_awprot),                         //                  .awprot
		.h2f_AWVALID              (hps_0_h2f_axi_master_awvalid),                        //                  .awvalid
		.h2f_AWREADY              (hps_0_h2f_axi_master_awready),                        //                  .awready
		.h2f_WID                  (hps_0_h2f_axi_master_wid),                            //                  .wid
		.h2f_WDATA                (hps_0_h2f_axi_master_wdata),                          //                  .wdata
		.h2f_WSTRB                (hps_0_h2f_axi_master_wstrb),                          //                  .wstrb
		.h2f_WLAST                (hps_0_h2f_axi_master_wlast),                          //                  .wlast
		.h2f_WVALID               (hps_0_h2f_axi_master_wvalid),                         //                  .wvalid
		.h2f_WREADY               (hps_0_h2f_axi_master_wready),                         //                  .wready
		.h2f_BID                  (hps_0_h2f_axi_master_bid),                            //                  .bid
		.h2f_BRESP                (hps_0_h2f_axi_master_bresp),                          //                  .bresp
		.h2f_BVALID               (hps_0_h2f_axi_master_bvalid),                         //                  .bvalid
		.h2f_BREADY               (hps_0_h2f_axi_master_bready),                         //                  .bready
		.h2f_ARID                 (hps_0_h2f_axi_master_arid),                           //                  .arid
		.h2f_ARADDR               (hps_0_h2f_axi_master_araddr),                         //                  .araddr
		.h2f_ARLEN                (hps_0_h2f_axi_master_arlen),                          //                  .arlen
		.h2f_ARSIZE               (hps_0_h2f_axi_master_arsize),                         //                  .arsize
		.h2f_ARBURST              (hps_0_h2f_axi_master_arburst),                        //                  .arburst
		.h2f_ARLOCK               (hps_0_h2f_axi_master_arlock),                         //                  .arlock
		.h2f_ARCACHE              (hps_0_h2f_axi_master_arcache),                        //                  .arcache
		.h2f_ARPROT               (hps_0_h2f_axi_master_arprot),                         //                  .arprot
		.h2f_ARVALID              (hps_0_h2f_axi_master_arvalid),                        //                  .arvalid
		.h2f_ARREADY              (hps_0_h2f_axi_master_arready),                        //                  .arready
		.h2f_RID                  (hps_0_h2f_axi_master_rid),                            //                  .rid
		.h2f_RDATA                (hps_0_h2f_axi_master_rdata),                          //                  .rdata
		.h2f_RRESP                (hps_0_h2f_axi_master_rresp),                          //                  .rresp
		.h2f_RLAST                (hps_0_h2f_axi_master_rlast),                          //                  .rlast
		.h2f_RVALID               (hps_0_h2f_axi_master_rvalid),                         //                  .rvalid
		.h2f_RREADY               (hps_0_h2f_axi_master_rready),                         //                  .rready
		.f2h_axi_clk              (clk_clk),                                             //     f2h_axi_clock.clk
		.f2h_AWID                 (hps_0_f2h_axi_slave_agent_altera_axi_master_awid),    //     f2h_axi_slave.awid
		.f2h_AWADDR               (hps_0_f2h_axi_slave_agent_altera_axi_master_awaddr),  //                  .awaddr
		.f2h_AWLEN                (hps_0_f2h_axi_slave_agent_altera_axi_master_awlen),   //                  .awlen
		.f2h_AWSIZE               (hps_0_f2h_axi_slave_agent_altera_axi_master_awsize),  //                  .awsize
		.f2h_AWBURST              (hps_0_f2h_axi_slave_agent_altera_axi_master_awburst), //                  .awburst
		.f2h_AWLOCK               (hps_0_f2h_axi_slave_agent_altera_axi_master_awlock),  //                  .awlock
		.f2h_AWCACHE              (hps_0_f2h_axi_slave_agent_altera_axi_master_awcache), //                  .awcache
		.f2h_AWPROT               (hps_0_f2h_axi_slave_agent_altera_axi_master_awprot),  //                  .awprot
		.f2h_AWVALID              (hps_0_f2h_axi_slave_agent_altera_axi_master_awvalid), //                  .awvalid
		.f2h_AWREADY              (hps_0_f2h_axi_slave_agent_altera_axi_master_awready), //                  .awready
		.f2h_AWUSER               (hps_0_f2h_axi_slave_agent_altera_axi_master_awuser),  //                  .awuser
		.f2h_WID                  (hps_0_f2h_axi_slave_agent_altera_axi_master_wid),     //                  .wid
		.f2h_WDATA                (hps_0_f2h_axi_slave_agent_altera_axi_master_wdata),   //                  .wdata
		.f2h_WSTRB                (hps_0_f2h_axi_slave_agent_altera_axi_master_wstrb),   //                  .wstrb
		.f2h_WLAST                (hps_0_f2h_axi_slave_agent_altera_axi_master_wlast),   //                  .wlast
		.f2h_WVALID               (hps_0_f2h_axi_slave_agent_altera_axi_master_wvalid),  //                  .wvalid
		.f2h_WREADY               (hps_0_f2h_axi_slave_agent_altera_axi_master_wready),  //                  .wready
		.f2h_BID                  (hps_0_f2h_axi_slave_agent_altera_axi_master_bid),     //                  .bid
		.f2h_BRESP                (hps_0_f2h_axi_slave_agent_altera_axi_master_bresp),   //                  .bresp
		.f2h_BVALID               (hps_0_f2h_axi_slave_agent_altera_axi_master_bvalid),  //                  .bvalid
		.f2h_BREADY               (hps_0_f2h_axi_slave_agent_altera_axi_master_bready),  //                  .bready
		.f2h_ARID                 (hps_0_f2h_axi_slave_agent_altera_axi_master_arid),    //                  .arid
		.f2h_ARADDR               (hps_0_f2h_axi_slave_agent_altera_axi_master_araddr),  //                  .araddr
		.f2h_ARLEN                (hps_0_f2h_axi_slave_agent_altera_axi_master_arlen),   //                  .arlen
		.f2h_ARSIZE               (hps_0_f2h_axi_slave_agent_altera_axi_master_arsize),  //                  .arsize
		.f2h_ARBURST              (hps_0_f2h_axi_slave_agent_altera_axi_master_arburst), //                  .arburst
		.f2h_ARLOCK               (hps_0_f2h_axi_slave_agent_altera_axi_master_arlock),  //                  .arlock
		.f2h_ARCACHE              (hps_0_f2h_axi_slave_agent_altera_axi_master_arcache), //                  .arcache
		.f2h_ARPROT               (hps_0_f2h_axi_slave_agent_altera_axi_master_arprot),  //                  .arprot
		.f2h_ARVALID              (hps_0_f2h_axi_slave_agent_altera_axi_master_arvalid), //                  .arvalid
		.f2h_ARREADY              (hps_0_f2h_axi_slave_agent_altera_axi_master_arready), //                  .arready
		.f2h_ARUSER               (hps_0_f2h_axi_slave_agent_altera_axi_master_aruser),  //                  .aruser
		.f2h_RID                  (hps_0_f2h_axi_slave_agent_altera_axi_master_rid),     //                  .rid
		.f2h_RDATA                (hps_0_f2h_axi_slave_agent_altera_axi_master_rdata),   //                  .rdata
		.f2h_RRESP                (hps_0_f2h_axi_slave_agent_altera_axi_master_rresp),   //                  .rresp
		.f2h_RLAST                (hps_0_f2h_axi_slave_agent_altera_axi_master_rlast),   //                  .rlast
		.f2h_RVALID               (hps_0_f2h_axi_slave_agent_altera_axi_master_rvalid),  //                  .rvalid
		.f2h_RREADY               (hps_0_f2h_axi_slave_agent_altera_axi_master_rready),  //                  .rready
		.h2f_lw_axi_clk           (clk_clk),                                             //  h2f_lw_axi_clock.clk
		.h2f_lw_AWID              (hps_0_h2f_lw_axi_master_awid),                        // h2f_lw_axi_master.awid
		.h2f_lw_AWADDR            (hps_0_h2f_lw_axi_master_awaddr),                      //                  .awaddr
		.h2f_lw_AWLEN             (hps_0_h2f_lw_axi_master_awlen),                       //                  .awlen
		.h2f_lw_AWSIZE            (hps_0_h2f_lw_axi_master_awsize),                      //                  .awsize
		.h2f_lw_AWBURST           (hps_0_h2f_lw_axi_master_awburst),                     //                  .awburst
		.h2f_lw_AWLOCK            (hps_0_h2f_lw_axi_master_awlock),                      //                  .awlock
		.h2f_lw_AWCACHE           (hps_0_h2f_lw_axi_master_awcache),                     //                  .awcache
		.h2f_lw_AWPROT            (hps_0_h2f_lw_axi_master_awprot),                      //                  .awprot
		.h2f_lw_AWVALID           (hps_0_h2f_lw_axi_master_awvalid),                     //                  .awvalid
		.h2f_lw_AWREADY           (hps_0_h2f_lw_axi_master_awready),                     //                  .awready
		.h2f_lw_WID               (hps_0_h2f_lw_axi_master_wid),                         //                  .wid
		.h2f_lw_WDATA             (hps_0_h2f_lw_axi_master_wdata),                       //                  .wdata
		.h2f_lw_WSTRB             (hps_0_h2f_lw_axi_master_wstrb),                       //                  .wstrb
		.h2f_lw_WLAST             (hps_0_h2f_lw_axi_master_wlast),                       //                  .wlast
		.h2f_lw_WVALID            (hps_0_h2f_lw_axi_master_wvalid),                      //                  .wvalid
		.h2f_lw_WREADY            (hps_0_h2f_lw_axi_master_wready),                      //                  .wready
		.h2f_lw_BID               (hps_0_h2f_lw_axi_master_bid),                         //                  .bid
		.h2f_lw_BRESP             (hps_0_h2f_lw_axi_master_bresp),                       //                  .bresp
		.h2f_lw_BVALID            (hps_0_h2f_lw_axi_master_bvalid),                      //                  .bvalid
		.h2f_lw_BREADY            (hps_0_h2f_lw_axi_master_bready),                      //                  .bready
		.h2f_lw_ARID              (hps_0_h2f_lw_axi_master_arid),                        //                  .arid
		.h2f_lw_ARADDR            (hps_0_h2f_lw_axi_master_araddr),                      //                  .araddr
		.h2f_lw_ARLEN             (hps_0_h2f_lw_axi_master_arlen),                       //                  .arlen
		.h2f_lw_ARSIZE            (hps_0_h2f_lw_axi_master_arsize),                      //                  .arsize
		.h2f_lw_ARBURST           (hps_0_h2f_lw_axi_master_arburst),                     //                  .arburst
		.h2f_lw_ARLOCK            (hps_0_h2f_lw_axi_master_arlock),                      //                  .arlock
		.h2f_lw_ARCACHE           (hps_0_h2f_lw_axi_master_arcache),                     //                  .arcache
		.h2f_lw_ARPROT            (hps_0_h2f_lw_axi_master_arprot),                      //                  .arprot
		.h2f_lw_ARVALID           (hps_0_h2f_lw_axi_master_arvalid),                     //                  .arvalid
		.h2f_lw_ARREADY           (hps_0_h2f_lw_axi_master_arready),                     //                  .arready
		.h2f_lw_RID               (hps_0_h2f_lw_axi_master_rid),                         //                  .rid
		.h2f_lw_RDATA             (hps_0_h2f_lw_axi_master_rdata),                       //                  .rdata
		.h2f_lw_RRESP             (hps_0_h2f_lw_axi_master_rresp),                       //                  .rresp
		.h2f_lw_RLAST             (hps_0_h2f_lw_axi_master_rlast),                       //                  .rlast
		.h2f_lw_RVALID            (hps_0_h2f_lw_axi_master_rvalid),                      //                  .rvalid
		.h2f_lw_RREADY            (hps_0_h2f_lw_axi_master_rready),                      //                  .rready
		.f2h_irq_p0               (hps_0_f2h_irq0_irq),                                  //          f2h_irq0.irq
		.f2h_irq_p1               (hps_0_f2h_irq1_irq)                                   //          f2h_irq1.irq
	);

	soc_system_master_secure #(
		.USE_PLI     (0),
		.PLI_PORT    (50000),
		.FIFO_DEPTHS (2)
	) master_secure (
		.clk_clk              (clk_clk),                            //          clk.clk
		.clk_reset_reset      (~reset_reset_n),                     //    clk_reset.reset
		.master_address       (master_secure_master_address),       //       master.address
		.master_readdata      (master_secure_master_readdata),      //             .readdata
		.master_read          (master_secure_master_read),          //             .read
		.master_write         (master_secure_master_write),         //             .write
		.master_writedata     (master_secure_master_writedata),     //             .writedata
		.master_waitrequest   (master_secure_master_waitrequest),   //             .waitrequest
		.master_readdatavalid (master_secure_master_readdatavalid), //             .readdatavalid
		.master_byteenable    (master_secure_master_byteenable),    //             .byteenable
		.master_reset_reset   ()                                    // master_reset.reset
	);

	soc_system_led_pio led_pio (
		.clk        (clk_clk),                                              //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                      //               reset.reset_n
		.address    (led_pio_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~led_pio_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (led_pio_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (led_pio_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (led_pio_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.out_port   (led_pio_external_connection_export)                    // external_connection.export
	);

	soc_system_dipsw_pio dipsw_pio (
		.clk        (clk_clk),                                                //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                        //               reset.reset_n
		.address    (dipsw_pio_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~dipsw_pio_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (dipsw_pio_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (dipsw_pio_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (dipsw_pio_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.in_port    (dipsw_pio_external_connection_export),                   // external_connection.export
		.irq        (irq_mapper_receiver2_irq)                                //                 irq.irq
	);

	soc_system_button_pio button_pio (
		.clk        (clk_clk),                                                 //                 clk.clk
		.reset_n    (~rst_controller_reset_out_reset),                         //               reset.reset_n
		.address    (button_pio_s1_translator_avalon_anti_slave_0_address),    //                  s1.address
		.write_n    (~button_pio_s1_translator_avalon_anti_slave_0_write),     //                    .write_n
		.writedata  (button_pio_s1_translator_avalon_anti_slave_0_writedata),  //                    .writedata
		.chipselect (button_pio_s1_translator_avalon_anti_slave_0_chipselect), //                    .chipselect
		.readdata   (button_pio_s1_translator_avalon_anti_slave_0_readdata),   //                    .readdata
		.in_port    (button_pio_external_connection_export),                   // external_connection.export
		.irq        (irq_mapper_receiver1_irq)                                 //                 irq.irq
	);

	soc_system_jtag_uart jtag_uart (
		.clk            (clk_clk),                                                                //               clk.clk
		.rst_n          (~rst_controller_reset_out_reset),                                        //             reset.reset_n
		.av_chipselect  (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect),  // avalon_jtag_slave.chipselect
		.av_address     (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_address),     //                  .address
		.av_read_n      (~jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read),       //                  .read_n
		.av_readdata    (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata),    //                  .readdata
		.av_write_n     (~jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write),      //                  .write_n
		.av_writedata   (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata),   //                  .writedata
		.av_waitrequest (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest), //                  .waitrequest
		.av_irq         (irq_mapper_receiver0_irq)                                                //               irq.irq
	);

	soc_system_pll_stream pll_stream (
		.refclk   (clk_clk),                        //  refclk.clk
		.rst      (rst_controller_reset_out_reset), //   reset.reset
		.outclk_0 (clock_bridge_148_5_out_clk_clk), // outclk0.clk
		.outclk_1 (pll_stream_outclk1_clk),         // outclk1.clk
		.locked   ()                                //  locked.export
	);

	soc_system_sdram sdram (
		.clk            (pll_sdram_outclk1_clk),                                 //   clk.clk
		.reset_n        (~rst_controller_001_reset_out_reset),                   // reset.reset_n
		.az_addr        (sdram_s1_translator_avalon_anti_slave_0_address),       //    s1.address
		.az_be_n        (~sdram_s1_translator_avalon_anti_slave_0_byteenable),   //      .byteenable_n
		.az_cs          (sdram_s1_translator_avalon_anti_slave_0_chipselect),    //      .chipselect
		.az_data        (sdram_s1_translator_avalon_anti_slave_0_writedata),     //      .writedata
		.az_rd_n        (~sdram_s1_translator_avalon_anti_slave_0_read),         //      .read_n
		.az_wr_n        (~sdram_s1_translator_avalon_anti_slave_0_write),        //      .write_n
		.za_data        (sdram_s1_translator_avalon_anti_slave_0_readdata),      //      .readdata
		.za_valid       (sdram_s1_translator_avalon_anti_slave_0_readdatavalid), //      .readdatavalid
		.za_waitrequest (sdram_s1_translator_avalon_anti_slave_0_waitrequest),   //      .waitrequest
		.zs_addr        (sdram_wire_addr),                                       //  wire.export
		.zs_ba          (sdram_wire_ba),                                         //      .export
		.zs_cas_n       (sdram_wire_cas_n),                                      //      .export
		.zs_cke         (sdram_wire_cke),                                        //      .export
		.zs_cs_n        (sdram_wire_cs_n),                                       //      .export
		.zs_dq          (sdram_wire_dq),                                         //      .export
		.zs_dqm         (sdram_wire_dqm),                                        //      .export
		.zs_ras_n       (sdram_wire_ras_n),                                      //      .export
		.zs_we_n        (sdram_wire_we_n)                                        //      .export
	);

	oc_i2c_master oc_i2c_master_0 (
		.wb_clk_i   (clk_clk),                                                                   //       clock_sink.clk
		.wb_rst_i   (rst_controller_reset_out_reset),                                            // clock_sink_reset.reset
		.wb_ack_o   (oc_i2c_master_0_avalon_slave_0_translator_avalon_anti_slave_0_waitrequest), //   avalon_slave_0.waitrequest_n
		.wb_adr_i   (oc_i2c_master_0_avalon_slave_0_translator_avalon_anti_slave_0_address),     //                 .address
		.wb_dat_i   (oc_i2c_master_0_avalon_slave_0_translator_avalon_anti_slave_0_writedata),   //                 .writedata
		.wb_dat_o   (oc_i2c_master_0_avalon_slave_0_translator_avalon_anti_slave_0_readdata),    //                 .readdata
		.wb_stb_i   (oc_i2c_master_0_avalon_slave_0_translator_avalon_anti_slave_0_chipselect),  //                 .chipselect
		.wb_we_i    (oc_i2c_master_0_avalon_slave_0_translator_avalon_anti_slave_0_write),       //                 .write
		.scl_pad_io (oc_i2c_master_0_conduit_start_scl_pad_io),                                  //    conduit_start.export
		.sda_pad_io (oc_i2c_master_0_conduit_start_sda_pad_io),                                  //                 .export
		.wb_inta_o  ()                                                                           // interrupt_sender.irq
	);

	soc_system_alt_vip_tpg_0 #(
		.CHANNELS_IN_PAR          (3),
		.CTRL_INTERFACE_DEPTH     (10),
		.PARAMETERISATION         ("<testPatternGeneratorParams><TPG_NAME>MyPatternGenerator</TPG_NAME><TPG_RUNTIME_CONTROL>0</TPG_RUNTIME_CONTROL><TPG_BPS>8</TPG_BPS><TPG_MAX_WIDTH>1280</TPG_MAX_WIDTH><TPG_MAX_HEIGHT>1024</TPG_MAX_HEIGHT><TPG_COLORSPACE>COLORSPACE_RGB</TPG_COLORSPACE><TPG_FORMAT>SAMPLE_444</TPG_FORMAT><TPG_INTERLACE>PROGRESSIVE_FRAMES</TPG_INTERLACE><TPG_PARALLEL_MODE>true</TPG_PARALLEL_MODE><TPG_PATTERN>TPG_PATTERN_UNIFORM</TPG_PATTERN><TPG_UNIFORM_VAL_C1>0</TPG_UNIFORM_VAL_C1><TPG_UNIFORM_VAL_C2>0</TPG_UNIFORM_VAL_C2><TPG_UNIFORM_VAL_C3>0</TPG_UNIFORM_VAL_C3></testPatternGeneratorParams>"),
		.AUTO_DEVICE_FAMILY       ("Cyclone V"),
		.AUTO_CONTROL_CLOCKS_SAME ("0")
	) alt_vip_tpg_0 (
		.clock              (pll_stream_outclk1_clk),             // clock.clk
		.reset              (rst_controller_002_reset_out_reset), // reset.reset
		.dout_ready         (alt_vip_tpg_0_dout_ready),           //  dout.ready
		.dout_valid         (alt_vip_tpg_0_dout_valid),           //      .valid
		.dout_data          (alt_vip_tpg_0_dout_data),            //      .data
		.dout_startofpacket (alt_vip_tpg_0_dout_startofpacket),   //      .startofpacket
		.dout_endofpacket   (alt_vip_tpg_0_dout_endofpacket)      //      .endofpacket
	);

	alt_vipvfr130_vfr #(
		.BITS_PER_PIXEL_PER_COLOR_PLANE (8),
		.NUMBER_OF_CHANNELS_IN_PARALLEL (3),
		.NUMBER_OF_CHANNELS_IN_SEQUENCE (1),
		.MAX_IMAGE_WIDTH                (640),
		.MAX_IMAGE_HEIGHT               (480),
		.MEM_PORT_WIDTH                 (32),
		.RMASTER_FIFO_DEPTH             (1024),
		.RMASTER_BURST_TARGET           (64),
		.CLOCKS_ARE_SEPARATE            (1)
	) alt_vip_vfr_0 (
		.clock                (pll_stream_outclk1_clk),                                              //             clock_reset.clk
		.reset                (rst_controller_002_reset_out_reset),                                  //       clock_reset_reset.reset
		.master_clock         (pll_sdram_outclk1_clk),                                               //            clock_master.clk
		.master_reset         (rst_controller_001_reset_out_reset),                                  //      clock_master_reset.reset
		.slave_address        (alt_vip_vfr_0_avalon_slave_translator_avalon_anti_slave_0_address),   //            avalon_slave.address
		.slave_write          (alt_vip_vfr_0_avalon_slave_translator_avalon_anti_slave_0_write),     //                        .write
		.slave_writedata      (alt_vip_vfr_0_avalon_slave_translator_avalon_anti_slave_0_writedata), //                        .writedata
		.slave_read           (alt_vip_vfr_0_avalon_slave_translator_avalon_anti_slave_0_read),      //                        .read
		.slave_readdata       (alt_vip_vfr_0_avalon_slave_translator_avalon_anti_slave_0_readdata),  //                        .readdata
		.slave_irq            (),                                                                    //        interrupt_sender.irq
		.dout_data            (alt_vip_vfr_0_avalon_streaming_source_data),                          // avalon_streaming_source.data
		.dout_valid           (alt_vip_vfr_0_avalon_streaming_source_valid),                         //                        .valid
		.dout_ready           (alt_vip_vfr_0_avalon_streaming_source_ready),                         //                        .ready
		.dout_startofpacket   (alt_vip_vfr_0_avalon_streaming_source_startofpacket),                 //                        .startofpacket
		.dout_endofpacket     (alt_vip_vfr_0_avalon_streaming_source_endofpacket),                   //                        .endofpacket
		.master_address       (alt_vip_vfr_0_avalon_master_address),                                 //           avalon_master.address
		.master_burstcount    (alt_vip_vfr_0_avalon_master_burstcount),                              //                        .burstcount
		.master_readdata      (alt_vip_vfr_0_avalon_master_readdata),                                //                        .readdata
		.master_read          (alt_vip_vfr_0_avalon_master_read),                                    //                        .read
		.master_readdatavalid (alt_vip_vfr_0_avalon_master_readdatavalid),                           //                        .readdatavalid
		.master_waitrequest   (alt_vip_vfr_0_avalon_master_waitrequest)                              //                        .waitrequest
	);

	soc_system_timing_adapter_0 timing_adapter_0 (
		.clk               (pll_stream_outclk1_clk),                //   clk.clk
		.reset_n           (~rst_controller_002_reset_out_reset),   // reset.reset_n
		.in_ready          (avalon_st_adapter_out_0_ready),         //    in.ready
		.in_valid          (avalon_st_adapter_out_0_valid),         //      .valid
		.in_data           (avalon_st_adapter_out_0_data),          //      .data
		.in_startofpacket  (avalon_st_adapter_out_0_startofpacket), //      .startofpacket
		.in_endofpacket    (avalon_st_adapter_out_0_endofpacket),   //      .endofpacket
		.out_ready         (timing_adapter_0_out_ready),            //   out.ready
		.out_valid         (timing_adapter_0_out_valid),            //      .valid
		.out_data          (timing_adapter_0_out_data),             //      .data
		.out_startofpacket (timing_adapter_0_out_startofpacket),    //      .startofpacket
		.out_endofpacket   (timing_adapter_0_out_endofpacket)       //      .endofpacket
	);

	soc_system_alt_vip_mix_0 #(
		.PARAMETERISATION         ("<mixerParams><MIX_NAME>mixer</MIX_NAME><MIX_ALPHA_ENABLED>false</MIX_ALPHA_ENABLED><MIX_ALPHA_BPS>8</MIX_ALPHA_BPS><MIX_CHANNELS_IN_SEQ>1</MIX_CHANNELS_IN_SEQ><MIX_CHANNELS_IN_PAR>3</MIX_CHANNELS_IN_PAR><MIX_BPS>8</MIX_BPS><MIX_NUM_LAYERS>3</MIX_NUM_LAYERS><MIX_RUNTIME_MAX_WIDTH>1280</MIX_RUNTIME_MAX_WIDTH><MIX_RUNTIME_MAX_HEIGHT>1024</MIX_RUNTIME_MAX_HEIGHT></mixerParams>"),
		.AUTO_DEVICE_FAMILY       ("Cyclone V"),
		.AUTO_CONTROL_CLOCKS_SAME ("2")
	) alt_vip_mix_0 (
		.clock                 (pll_stream_outclk1_clk),                                          //   clock.clk
		.reset                 (rst_controller_002_reset_out_reset),                              //   reset.reset
		.din_0_ready           (alt_vip_tpg_0_dout_ready),                                        //   din_0.ready
		.din_0_valid           (alt_vip_tpg_0_dout_valid),                                        //        .valid
		.din_0_data            (alt_vip_tpg_0_dout_data),                                         //        .data
		.din_0_startofpacket   (alt_vip_tpg_0_dout_startofpacket),                                //        .startofpacket
		.din_0_endofpacket     (alt_vip_tpg_0_dout_endofpacket),                                  //        .endofpacket
		.din_1_ready           (timing_adapter_0_out_ready),                                      //   din_1.ready
		.din_1_valid           (timing_adapter_0_out_valid),                                      //        .valid
		.din_1_data            (timing_adapter_0_out_data),                                       //        .data
		.din_1_startofpacket   (timing_adapter_0_out_startofpacket),                              //        .startofpacket
		.din_1_endofpacket     (timing_adapter_0_out_endofpacket),                                //        .endofpacket
		.din_2_ready           (alt_vip_vfr_0_avalon_streaming_source_ready),                     //   din_2.ready
		.din_2_valid           (alt_vip_vfr_0_avalon_streaming_source_valid),                     //        .valid
		.din_2_data            (alt_vip_vfr_0_avalon_streaming_source_data),                      //        .data
		.din_2_startofpacket   (alt_vip_vfr_0_avalon_streaming_source_startofpacket),             //        .startofpacket
		.din_2_endofpacket     (alt_vip_vfr_0_avalon_streaming_source_endofpacket),               //        .endofpacket
		.dout_ready            (alt_vip_mix_0_dout_ready),                                        //    dout.ready
		.dout_valid            (alt_vip_mix_0_dout_valid),                                        //        .valid
		.dout_data             (alt_vip_mix_0_dout_data),                                         //        .data
		.dout_startofpacket    (alt_vip_mix_0_dout_startofpacket),                                //        .startofpacket
		.dout_endofpacket      (alt_vip_mix_0_dout_endofpacket),                                  //        .endofpacket
		.control_av_chipselect (alt_vip_mix_0_control_translator_avalon_anti_slave_0_chipselect), // control.chipselect
		.control_av_write      (alt_vip_mix_0_control_translator_avalon_anti_slave_0_write),      //        .write
		.control_av_address    (alt_vip_mix_0_control_translator_avalon_anti_slave_0_address),    //        .address
		.control_av_writedata  (alt_vip_mix_0_control_translator_avalon_anti_slave_0_writedata),  //        .writedata
		.control_av_readdata   (alt_vip_mix_0_control_translator_avalon_anti_slave_0_readdata)    //        .readdata
	);

	alt_vipitc130_IS2Vid #(
		.NUMBER_OF_COLOUR_PLANES       (3),
		.COLOUR_PLANES_ARE_IN_PARALLEL (1),
		.BPS                           (8),
		.INTERLACED                    (0),
		.H_ACTIVE_PIXELS               (1280),
		.V_ACTIVE_LINES                (1024),
		.ACCEPT_COLOURS_IN_SEQ         (0),
		.FIFO_DEPTH                    (1280),
		.CLOCKS_ARE_SAME               (0),
		.USE_CONTROL                   (0),
		.NO_OF_MODES                   (1),
		.THRESHOLD                     (1279),
		.STD_WIDTH                     (1),
		.GENERATE_SYNC                 (0),
		.USE_EMBEDDED_SYNCS            (0),
		.AP_LINE                       (0),
		.V_BLANK                       (0),
		.H_BLANK                       (0),
		.H_SYNC_LENGTH                 (112),
		.H_FRONT_PORCH                 (48),
		.H_BACK_PORCH                  (248),
		.V_SYNC_LENGTH                 (3),
		.V_FRONT_PORCH                 (1),
		.V_BACK_PORCH                  (38),
		.F_RISING_EDGE                 (0),
		.F_FALLING_EDGE                (0),
		.FIELD0_V_RISING_EDGE          (0),
		.FIELD0_V_BLANK                (0),
		.FIELD0_V_SYNC_LENGTH          (0),
		.FIELD0_V_FRONT_PORCH          (0),
		.FIELD0_V_BACK_PORCH           (0),
		.ANC_LINE                      (0),
		.FIELD0_ANC_LINE               (0)
	) alt_vip_itc_0 (
		.is_clk        (pll_stream_outclk1_clk),                    //       is_clk_rst.clk
		.rst           (rst_controller_002_reset_out_reset),        // is_clk_rst_reset.reset
		.is_data       (alt_vip_mix_0_dout_data),                   //              din.data
		.is_valid      (alt_vip_mix_0_dout_valid),                  //                 .valid
		.is_ready      (alt_vip_mix_0_dout_ready),                  //                 .ready
		.is_sop        (alt_vip_mix_0_dout_startofpacket),          //                 .startofpacket
		.is_eop        (alt_vip_mix_0_dout_endofpacket),            //                 .endofpacket
		.vid_clk       (alt_vip_itc_0_clocked_video_vid_clk),       //    clocked_video.export
		.vid_data      (alt_vip_itc_0_clocked_video_vid_data),      //                 .export
		.underflow     (alt_vip_itc_0_clocked_video_underflow),     //                 .export
		.vid_datavalid (alt_vip_itc_0_clocked_video_vid_datavalid), //                 .export
		.vid_v_sync    (alt_vip_itc_0_clocked_video_vid_v_sync),    //                 .export
		.vid_h_sync    (alt_vip_itc_0_clocked_video_vid_h_sync),    //                 .export
		.vid_f         (alt_vip_itc_0_clocked_video_vid_f),         //                 .export
		.vid_h         (alt_vip_itc_0_clocked_video_vid_h),         //                 .export
		.vid_v         (alt_vip_itc_0_clocked_video_vid_v)          //                 .export
	);

	soc_system_pll_sdram pll_sdram (
		.refclk   (clk_clk),                        //  refclk.clk
		.rst      (rst_controller_reset_out_reset), //   reset.reset
		.outclk_0 (sdram_clk_clk),                  // outclk0.clk
		.outclk_1 (pll_sdram_outclk1_clk),          // outclk1.clk
		.locked   ()                                //  locked.export
	);

	soc_system_pll_audio pll_audio (
		.refclk   (clk_clk),                        //  refclk.clk
		.rst      (rst_controller_reset_out_reset), //   reset.reset
		.outclk_0 (pll_audio_outclk0_clk),          // outclk0.clk
		.locked   ()                                //  locked.export
	);

	log_generator #(
		.BACK_COLOR        (26'b00000000000000000000000001),
		.FRONT_COLOR       (26'b00111111111111111111111111),
		.MIF_FILE_LOCATION ("./log.mif"),
		.LOG_WIDTH         (1024),
		.LOG_HEIGHT        (249)
	) log_generate_0 (
		.reset      (rst_controller_002_reset_out_reset), //      reset.reset
		.clock      (pll_stream_outclk1_clk),             // clock_sink.clk
		.dout_ready (log_generate_0_dout_ready),          //       dout.ready
		.dout_valid (log_generate_0_dout_valid),          //           .valid
		.dout_data  (log_generate_0_dout_data),           //           .data
		.dout_sop   (log_generate_0_dout_startofpacket),  //           .startofpacket
		.dout_eop   (log_generate_0_dout_endofpacket),    //           .endofpacket
		.dout_empty (log_generate_0_dout_empty)           //           .empty
	);

	AUDIO_IF audio_if_0 (
		.avs_s1_address       (audio_if_0_avalon_slave_translator_avalon_anti_slave_0_address),   //     avalon_slave.address
		.avs_s1_read          (audio_if_0_avalon_slave_translator_avalon_anti_slave_0_read),      //                 .read
		.avs_s1_readdata      (audio_if_0_avalon_slave_translator_avalon_anti_slave_0_readdata),  //                 .readdata
		.avs_s1_write         (audio_if_0_avalon_slave_translator_avalon_anti_slave_0_write),     //                 .write
		.avs_s1_writedata     (audio_if_0_avalon_slave_translator_avalon_anti_slave_0_writedata), //                 .writedata
		.avs_s1_clk           (pll_audio_outclk0_clk),                                            //       clock_sink.clk
		.avs_s1_reset         (rst_controller_003_reset_out_reset),                               // clock_sink_reset.reset
		.avs_s1_export_XCK    (audio_if_0_conduit_end_XCK),                                       //      conduit_end.export
		.avs_s1_export_ADCDAT (audio_if_0_conduit_end_ADCDAT),                                    //                 .export
		.avs_s1_export_ADCLRC (audio_if_0_conduit_end_ADCLRC),                                    //                 .export
		.avs_s1_export_DACDAT (audio_if_0_conduit_end_DACDAT),                                    //                 .export
		.avs_s1_export_DACLRC (audio_if_0_conduit_end_DACLRC),                                    //                 .export
		.avs_s1_export_BCLK   (audio_if_0_conduit_end_BCLK)                                       //                 .export
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (32),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (1),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (3),
		.USE_READ                    (1),
		.USE_WRITE                   (1),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (0),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.USE_READRESPONSE            (0),
		.USE_WRITERESPONSE           (0),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (0),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) master_secure_master_translator (
		.clk                      (clk_clk),                                                                 //                       clk.clk
		.reset                    (rst_controller_reset_out_reset),                                          //                     reset.reset
		.uav_address              (master_secure_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount           (master_secure_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read                 (master_secure_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write                (master_secure_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest          (master_secure_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid        (master_secure_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable           (master_secure_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata             (master_secure_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata            (master_secure_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock                 (master_secure_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess          (master_secure_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address               (master_secure_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest           (master_secure_master_waitrequest),                                        //                          .waitrequest
		.av_byteenable            (master_secure_master_byteenable),                                         //                          .byteenable
		.av_read                  (master_secure_master_read),                                               //                          .read
		.av_readdata              (master_secure_master_readdata),                                           //                          .readdata
		.av_readdatavalid         (master_secure_master_readdatavalid),                                      //                          .readdatavalid
		.av_write                 (master_secure_master_write),                                              //                          .write
		.av_writedata             (master_secure_master_writedata),                                          //                          .writedata
		.av_burstcount            (1'b1),                                                                    //               (terminated)
		.av_beginbursttransfer    (1'b0),                                                                    //               (terminated)
		.av_begintransfer         (1'b0),                                                                    //               (terminated)
		.av_chipselect            (1'b0),                                                                    //               (terminated)
		.av_lock                  (1'b0),                                                                    //               (terminated)
		.av_debugaccess           (1'b0),                                                                    //               (terminated)
		.uav_clken                (),                                                                        //               (terminated)
		.av_clken                 (1'b1),                                                                    //               (terminated)
		.uav_response             (2'b00),                                                                   //               (terminated)
		.av_response              (),                                                                        //               (terminated)
		.uav_writeresponserequest (),                                                                        //               (terminated)
		.uav_writeresponsevalid   (1'b0),                                                                    //               (terminated)
		.av_writeresponserequest  (1'b0),                                                                    //               (terminated)
		.av_writeresponsevalid    ()                                                                         //               (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (21),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) led_pio_s1_translator (
		.clk                      (clk_clk),                                                               //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                        //                    reset.reset
		.uav_address              (led_pio_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (led_pio_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (led_pio_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (led_pio_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (led_pio_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (led_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (led_pio_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (led_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (led_pio_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (led_pio_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (led_pio_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (led_pio_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (led_pio_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (led_pio_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (led_pio_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (led_pio_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                      //              (terminated)
		.av_begintransfer         (),                                                                      //              (terminated)
		.av_beginbursttransfer    (),                                                                      //              (terminated)
		.av_burstcount            (),                                                                      //              (terminated)
		.av_byteenable            (),                                                                      //              (terminated)
		.av_readdatavalid         (1'b0),                                                                  //              (terminated)
		.av_waitrequest           (1'b0),                                                                  //              (terminated)
		.av_writebyteenable       (),                                                                      //              (terminated)
		.av_lock                  (),                                                                      //              (terminated)
		.av_clken                 (),                                                                      //              (terminated)
		.uav_clken                (1'b0),                                                                  //              (terminated)
		.av_debugaccess           (),                                                                      //              (terminated)
		.av_outputenable          (),                                                                      //              (terminated)
		.uav_response             (),                                                                      //              (terminated)
		.av_response              (2'b00),                                                                 //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                  //              (terminated)
		.uav_writeresponsevalid   (),                                                                      //              (terminated)
		.av_writeresponserequest  (),                                                                      //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                   //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (21),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) dipsw_pio_s1_translator (
		.clk                      (clk_clk),                                                                 //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                          //                    reset.reset
		.uav_address              (dipsw_pio_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (dipsw_pio_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (dipsw_pio_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (dipsw_pio_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (dipsw_pio_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (dipsw_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (dipsw_pio_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (dipsw_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (dipsw_pio_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (dipsw_pio_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (dipsw_pio_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (dipsw_pio_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (dipsw_pio_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (dipsw_pio_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (dipsw_pio_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (dipsw_pio_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                        //              (terminated)
		.av_begintransfer         (),                                                                        //              (terminated)
		.av_beginbursttransfer    (),                                                                        //              (terminated)
		.av_burstcount            (),                                                                        //              (terminated)
		.av_byteenable            (),                                                                        //              (terminated)
		.av_readdatavalid         (1'b0),                                                                    //              (terminated)
		.av_waitrequest           (1'b0),                                                                    //              (terminated)
		.av_writebyteenable       (),                                                                        //              (terminated)
		.av_lock                  (),                                                                        //              (terminated)
		.av_clken                 (),                                                                        //              (terminated)
		.uav_clken                (1'b0),                                                                    //              (terminated)
		.av_debugaccess           (),                                                                        //              (terminated)
		.av_outputenable          (),                                                                        //              (terminated)
		.uav_response             (),                                                                        //              (terminated)
		.av_response              (2'b00),                                                                   //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                    //              (terminated)
		.uav_writeresponsevalid   (),                                                                        //              (terminated)
		.av_writeresponserequest  (),                                                                        //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                     //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (2),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (21),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) button_pio_s1_translator (
		.clk                      (clk_clk),                                                                  //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                           //                    reset.reset
		.uav_address              (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (button_pio_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (button_pio_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (button_pio_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (button_pio_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (button_pio_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                         //              (terminated)
		.av_begintransfer         (),                                                                         //              (terminated)
		.av_beginbursttransfer    (),                                                                         //              (terminated)
		.av_burstcount            (),                                                                         //              (terminated)
		.av_byteenable            (),                                                                         //              (terminated)
		.av_readdatavalid         (1'b0),                                                                     //              (terminated)
		.av_waitrequest           (1'b0),                                                                     //              (terminated)
		.av_writebyteenable       (),                                                                         //              (terminated)
		.av_lock                  (),                                                                         //              (terminated)
		.av_clken                 (),                                                                         //              (terminated)
		.uav_clken                (1'b0),                                                                     //              (terminated)
		.av_debugaccess           (),                                                                         //              (terminated)
		.av_outputenable          (),                                                                         //              (terminated)
		.uav_response             (),                                                                         //              (terminated)
		.av_response              (2'b00),                                                                    //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                     //              (terminated)
		.uav_writeresponsevalid   (),                                                                         //              (terminated)
		.av_writeresponserequest  (),                                                                         //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                      //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (1),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (21),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) jtag_uart_avalon_jtag_slave_translator (
		.clk                      (clk_clk),                                                                                //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                         //                    reset.reset
		.uav_address              (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest           (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_chipselect            (jtag_uart_avalon_jtag_slave_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer         (),                                                                                       //              (terminated)
		.av_beginbursttransfer    (),                                                                                       //              (terminated)
		.av_burstcount            (),                                                                                       //              (terminated)
		.av_byteenable            (),                                                                                       //              (terminated)
		.av_readdatavalid         (1'b0),                                                                                   //              (terminated)
		.av_writebyteenable       (),                                                                                       //              (terminated)
		.av_lock                  (),                                                                                       //              (terminated)
		.av_clken                 (),                                                                                       //              (terminated)
		.uav_clken                (1'b0),                                                                                   //              (terminated)
		.av_debugaccess           (),                                                                                       //              (terminated)
		.av_outputenable          (),                                                                                       //              (terminated)
		.uav_response             (),                                                                                       //              (terminated)
		.av_response              (2'b00),                                                                                  //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                   //              (terminated)
		.uav_writeresponsevalid   (),                                                                                       //              (terminated)
		.av_writeresponserequest  (),                                                                                       //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                    //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (4),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (21),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) oc_i2c_master_0_avalon_slave_0_translator (
		.clk                      (clk_clk),                                                                                   //                      clk.clk
		.reset                    (rst_controller_reset_out_reset),                                                            //                    reset.reset
		.uav_address              (oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (oc_i2c_master_0_avalon_slave_0_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (oc_i2c_master_0_avalon_slave_0_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (oc_i2c_master_0_avalon_slave_0_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (oc_i2c_master_0_avalon_slave_0_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_waitrequest           (~oc_i2c_master_0_avalon_slave_0_translator_avalon_anti_slave_0_waitrequest),                //                         .waitrequest
		.av_chipselect            (oc_i2c_master_0_avalon_slave_0_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                                          //              (terminated)
		.av_begintransfer         (),                                                                                          //              (terminated)
		.av_beginbursttransfer    (),                                                                                          //              (terminated)
		.av_burstcount            (),                                                                                          //              (terminated)
		.av_byteenable            (),                                                                                          //              (terminated)
		.av_readdatavalid         (1'b0),                                                                                      //              (terminated)
		.av_writebyteenable       (),                                                                                          //              (terminated)
		.av_lock                  (),                                                                                          //              (terminated)
		.av_clken                 (),                                                                                          //              (terminated)
		.uav_clken                (1'b0),                                                                                      //              (terminated)
		.av_debugaccess           (),                                                                                          //              (terminated)
		.av_outputenable          (),                                                                                          //              (terminated)
		.uav_response             (),                                                                                          //              (terminated)
		.av_response              (2'b00),                                                                                     //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                      //              (terminated)
		.uav_writeresponsevalid   (),                                                                                          //              (terminated)
		.av_writeresponserequest  (),                                                                                          //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                       //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (6),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (21),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (2),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) alt_vip_mix_0_control_translator (
		.clk                      (pll_stream_outclk1_clk),                                                           //                      clk.clk
		.reset                    (rst_controller_002_reset_out_reset),                                               //                    reset.reset
		.uav_address              (alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (alt_vip_mix_0_control_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (alt_vip_mix_0_control_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_readdata              (alt_vip_mix_0_control_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (alt_vip_mix_0_control_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_chipselect            (alt_vip_mix_0_control_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_read                  (),                                                                                 //              (terminated)
		.av_begintransfer         (),                                                                                 //              (terminated)
		.av_beginbursttransfer    (),                                                                                 //              (terminated)
		.av_burstcount            (),                                                                                 //              (terminated)
		.av_byteenable            (),                                                                                 //              (terminated)
		.av_readdatavalid         (1'b0),                                                                             //              (terminated)
		.av_waitrequest           (1'b0),                                                                             //              (terminated)
		.av_writebyteenable       (),                                                                                 //              (terminated)
		.av_lock                  (),                                                                                 //              (terminated)
		.av_clken                 (),                                                                                 //              (terminated)
		.uav_clken                (1'b0),                                                                             //              (terminated)
		.av_debugaccess           (),                                                                                 //              (terminated)
		.av_outputenable          (),                                                                                 //              (terminated)
		.uav_response             (),                                                                                 //              (terminated)
		.av_response              (2'b00),                                                                            //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                             //              (terminated)
		.uav_writeresponsevalid   (),                                                                                 //              (terminated)
		.av_writeresponserequest  (),                                                                                 //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                              //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (5),
		.AV_DATA_W                      (32),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (21),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (1),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) alt_vip_vfr_0_avalon_slave_translator (
		.clk                      (pll_stream_outclk1_clk),                                                                //                      clk.clk
		.reset                    (rst_controller_002_reset_out_reset),                                                    //                    reset.reset
		.uav_address              (alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (alt_vip_vfr_0_avalon_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (alt_vip_vfr_0_avalon_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (alt_vip_vfr_0_avalon_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (alt_vip_vfr_0_avalon_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (alt_vip_vfr_0_avalon_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_begintransfer         (),                                                                                      //              (terminated)
		.av_beginbursttransfer    (),                                                                                      //              (terminated)
		.av_burstcount            (),                                                                                      //              (terminated)
		.av_byteenable            (),                                                                                      //              (terminated)
		.av_readdatavalid         (1'b0),                                                                                  //              (terminated)
		.av_waitrequest           (1'b0),                                                                                  //              (terminated)
		.av_writebyteenable       (),                                                                                      //              (terminated)
		.av_lock                  (),                                                                                      //              (terminated)
		.av_chipselect            (),                                                                                      //              (terminated)
		.av_clken                 (),                                                                                      //              (terminated)
		.uav_clken                (1'b0),                                                                                  //              (terminated)
		.av_debugaccess           (),                                                                                      //              (terminated)
		.av_outputenable          (),                                                                                      //              (terminated)
		.uav_response             (),                                                                                      //              (terminated)
		.av_response              (2'b00),                                                                                 //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                                  //              (terminated)
		.uav_writeresponsevalid   (),                                                                                      //              (terminated)
		.av_writeresponserequest  (),                                                                                      //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                   //              (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (3),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (32),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (1),
		.UAV_BYTEENABLE_W               (4),
		.UAV_ADDRESS_W                  (21),
		.UAV_BURSTCOUNT_W               (3),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (0),
		.USE_WAITREQUEST                (0),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (4),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (0),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) audio_if_0_avalon_slave_translator (
		.clk                      (pll_audio_outclk0_clk),                                                              //                      clk.clk
		.reset                    (rst_controller_003_reset_out_reset),                                                 //                    reset.reset
		.uav_address              (audio_if_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (audio_if_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (audio_if_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (audio_if_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (audio_if_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (audio_if_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (audio_if_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (audio_if_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (audio_if_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (audio_if_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (audio_if_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (audio_if_0_avalon_slave_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (audio_if_0_avalon_slave_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (audio_if_0_avalon_slave_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (audio_if_0_avalon_slave_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (audio_if_0_avalon_slave_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_begintransfer         (),                                                                                   //              (terminated)
		.av_beginbursttransfer    (),                                                                                   //              (terminated)
		.av_burstcount            (),                                                                                   //              (terminated)
		.av_byteenable            (),                                                                                   //              (terminated)
		.av_readdatavalid         (1'b0),                                                                               //              (terminated)
		.av_waitrequest           (1'b0),                                                                               //              (terminated)
		.av_writebyteenable       (),                                                                                   //              (terminated)
		.av_lock                  (),                                                                                   //              (terminated)
		.av_chipselect            (),                                                                                   //              (terminated)
		.av_clken                 (),                                                                                   //              (terminated)
		.uav_clken                (1'b0),                                                                               //              (terminated)
		.av_debugaccess           (),                                                                                   //              (terminated)
		.av_outputenable          (),                                                                                   //              (terminated)
		.uav_response             (),                                                                                   //              (terminated)
		.av_response              (2'b00),                                                                              //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                               //              (terminated)
		.uav_writeresponsevalid   (),                                                                                   //              (terminated)
		.av_writeresponserequest  (),                                                                                   //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                                //              (terminated)
	);

	altera_merlin_master_translator #(
		.AV_ADDRESS_W                (32),
		.AV_DATA_W                   (32),
		.AV_BURSTCOUNT_W             (7),
		.AV_BYTEENABLE_W             (4),
		.UAV_ADDRESS_W               (32),
		.UAV_BURSTCOUNT_W            (9),
		.USE_READ                    (1),
		.USE_WRITE                   (0),
		.USE_BEGINBURSTTRANSFER      (0),
		.USE_BEGINTRANSFER           (0),
		.USE_CHIPSELECT              (0),
		.USE_BURSTCOUNT              (1),
		.USE_READDATAVALID           (1),
		.USE_WAITREQUEST             (1),
		.USE_READRESPONSE            (0),
		.USE_WRITERESPONSE           (0),
		.AV_SYMBOLS_PER_WORD         (4),
		.AV_ADDRESS_SYMBOLS          (1),
		.AV_BURSTCOUNT_SYMBOLS       (0),
		.AV_CONSTANT_BURST_BEHAVIOR  (1),
		.UAV_CONSTANT_BURST_BEHAVIOR (0),
		.AV_LINEWRAPBURSTS           (0),
		.AV_REGISTERINCOMINGSIGNALS  (0)
	) alt_vip_vfr_0_avalon_master_translator (
		.clk                      (pll_sdram_outclk1_clk),                                                          //                       clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                             //                     reset.reset
		.uav_address              (alt_vip_vfr_0_avalon_master_translator_avalon_universal_master_0_address),       // avalon_universal_master_0.address
		.uav_burstcount           (alt_vip_vfr_0_avalon_master_translator_avalon_universal_master_0_burstcount),    //                          .burstcount
		.uav_read                 (alt_vip_vfr_0_avalon_master_translator_avalon_universal_master_0_read),          //                          .read
		.uav_write                (alt_vip_vfr_0_avalon_master_translator_avalon_universal_master_0_write),         //                          .write
		.uav_waitrequest          (alt_vip_vfr_0_avalon_master_translator_avalon_universal_master_0_waitrequest),   //                          .waitrequest
		.uav_readdatavalid        (alt_vip_vfr_0_avalon_master_translator_avalon_universal_master_0_readdatavalid), //                          .readdatavalid
		.uav_byteenable           (alt_vip_vfr_0_avalon_master_translator_avalon_universal_master_0_byteenable),    //                          .byteenable
		.uav_readdata             (alt_vip_vfr_0_avalon_master_translator_avalon_universal_master_0_readdata),      //                          .readdata
		.uav_writedata            (alt_vip_vfr_0_avalon_master_translator_avalon_universal_master_0_writedata),     //                          .writedata
		.uav_lock                 (alt_vip_vfr_0_avalon_master_translator_avalon_universal_master_0_lock),          //                          .lock
		.uav_debugaccess          (alt_vip_vfr_0_avalon_master_translator_avalon_universal_master_0_debugaccess),   //                          .debugaccess
		.av_address               (alt_vip_vfr_0_avalon_master_address),                                            //      avalon_anti_master_0.address
		.av_waitrequest           (alt_vip_vfr_0_avalon_master_waitrequest),                                        //                          .waitrequest
		.av_burstcount            (alt_vip_vfr_0_avalon_master_burstcount),                                         //                          .burstcount
		.av_read                  (alt_vip_vfr_0_avalon_master_read),                                               //                          .read
		.av_readdata              (alt_vip_vfr_0_avalon_master_readdata),                                           //                          .readdata
		.av_readdatavalid         (alt_vip_vfr_0_avalon_master_readdatavalid),                                      //                          .readdatavalid
		.av_byteenable            (4'b1111),                                                                        //               (terminated)
		.av_beginbursttransfer    (1'b0),                                                                           //               (terminated)
		.av_begintransfer         (1'b0),                                                                           //               (terminated)
		.av_chipselect            (1'b0),                                                                           //               (terminated)
		.av_write                 (1'b0),                                                                           //               (terminated)
		.av_writedata             (32'b00000000000000000000000000000000),                                           //               (terminated)
		.av_lock                  (1'b0),                                                                           //               (terminated)
		.av_debugaccess           (1'b0),                                                                           //               (terminated)
		.uav_clken                (),                                                                               //               (terminated)
		.av_clken                 (1'b1),                                                                           //               (terminated)
		.uav_response             (2'b00),                                                                          //               (terminated)
		.av_response              (),                                                                               //               (terminated)
		.uav_writeresponserequest (),                                                                               //               (terminated)
		.uav_writeresponsevalid   (1'b0),                                                                           //               (terminated)
		.av_writeresponserequest  (1'b0),                                                                           //               (terminated)
		.av_writeresponsevalid    ()                                                                                //               (terminated)
	);

	altera_merlin_slave_translator #(
		.AV_ADDRESS_W                   (25),
		.AV_DATA_W                      (16),
		.UAV_DATA_W                     (16),
		.AV_BURSTCOUNT_W                (1),
		.AV_BYTEENABLE_W                (2),
		.UAV_BYTEENABLE_W               (2),
		.UAV_ADDRESS_W                  (32),
		.UAV_BURSTCOUNT_W               (2),
		.AV_READLATENCY                 (0),
		.USE_READDATAVALID              (1),
		.USE_WAITREQUEST                (1),
		.USE_UAV_CLKEN                  (0),
		.USE_READRESPONSE               (0),
		.USE_WRITERESPONSE              (0),
		.AV_SYMBOLS_PER_WORD            (2),
		.AV_ADDRESS_SYMBOLS             (0),
		.AV_BURSTCOUNT_SYMBOLS          (0),
		.AV_CONSTANT_BURST_BEHAVIOR     (0),
		.UAV_CONSTANT_BURST_BEHAVIOR    (0),
		.AV_REQUIRE_UNALIGNED_ADDRESSES (0),
		.CHIPSELECT_THROUGH_READLATENCY (0),
		.AV_READ_WAIT_CYCLES            (1),
		.AV_WRITE_WAIT_CYCLES           (0),
		.AV_SETUP_WAIT_CYCLES           (0),
		.AV_DATA_HOLD_CYCLES            (0)
	) sdram_s1_translator (
		.clk                      (pll_sdram_outclk1_clk),                                               //                      clk.clk
		.reset                    (rst_controller_001_reset_out_reset),                                  //                    reset.reset
		.uav_address              (sdram_s1_translator_avalon_universal_slave_0_agent_m0_address),       // avalon_universal_slave_0.address
		.uav_burstcount           (sdram_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),    //                         .burstcount
		.uav_read                 (sdram_s1_translator_avalon_universal_slave_0_agent_m0_read),          //                         .read
		.uav_write                (sdram_s1_translator_avalon_universal_slave_0_agent_m0_write),         //                         .write
		.uav_waitrequest          (sdram_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),   //                         .waitrequest
		.uav_readdatavalid        (sdram_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid), //                         .readdatavalid
		.uav_byteenable           (sdram_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),    //                         .byteenable
		.uav_readdata             (sdram_s1_translator_avalon_universal_slave_0_agent_m0_readdata),      //                         .readdata
		.uav_writedata            (sdram_s1_translator_avalon_universal_slave_0_agent_m0_writedata),     //                         .writedata
		.uav_lock                 (sdram_s1_translator_avalon_universal_slave_0_agent_m0_lock),          //                         .lock
		.uav_debugaccess          (sdram_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),   //                         .debugaccess
		.av_address               (sdram_s1_translator_avalon_anti_slave_0_address),                     //      avalon_anti_slave_0.address
		.av_write                 (sdram_s1_translator_avalon_anti_slave_0_write),                       //                         .write
		.av_read                  (sdram_s1_translator_avalon_anti_slave_0_read),                        //                         .read
		.av_readdata              (sdram_s1_translator_avalon_anti_slave_0_readdata),                    //                         .readdata
		.av_writedata             (sdram_s1_translator_avalon_anti_slave_0_writedata),                   //                         .writedata
		.av_byteenable            (sdram_s1_translator_avalon_anti_slave_0_byteenable),                  //                         .byteenable
		.av_readdatavalid         (sdram_s1_translator_avalon_anti_slave_0_readdatavalid),               //                         .readdatavalid
		.av_waitrequest           (sdram_s1_translator_avalon_anti_slave_0_waitrequest),                 //                         .waitrequest
		.av_chipselect            (sdram_s1_translator_avalon_anti_slave_0_chipselect),                  //                         .chipselect
		.av_begintransfer         (),                                                                    //              (terminated)
		.av_beginbursttransfer    (),                                                                    //              (terminated)
		.av_burstcount            (),                                                                    //              (terminated)
		.av_writebyteenable       (),                                                                    //              (terminated)
		.av_lock                  (),                                                                    //              (terminated)
		.av_clken                 (),                                                                    //              (terminated)
		.uav_clken                (1'b0),                                                                //              (terminated)
		.av_debugaccess           (),                                                                    //              (terminated)
		.av_outputenable          (),                                                                    //              (terminated)
		.uav_response             (),                                                                    //              (terminated)
		.av_response              (2'b00),                                                               //              (terminated)
		.uav_writeresponserequest (1'b0),                                                                //              (terminated)
		.uav_writeresponsevalid   (),                                                                    //              (terminated)
		.av_writeresponserequest  (),                                                                    //              (terminated)
		.av_writeresponsevalid    (1'b0)                                                                 //              (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (108),
		.PKT_PROTECTION_L          (106),
		.PKT_BEGIN_BURST           (101),
		.PKT_BURSTWRAP_H           (89),
		.PKT_BURSTWRAP_L           (82),
		.PKT_BURST_SIZE_H          (92),
		.PKT_BURST_SIZE_L          (90),
		.PKT_BURST_TYPE_H          (94),
		.PKT_BURST_TYPE_L          (93),
		.PKT_BYTE_CNT_H            (81),
		.PKT_BYTE_CNT_L            (74),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_TRANS_EXCLUSIVE       (73),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (103),
		.PKT_SRC_ID_L              (103),
		.PKT_DEST_ID_H             (104),
		.PKT_DEST_ID_L             (104),
		.PKT_THREAD_ID_H           (105),
		.PKT_THREAD_ID_L           (105),
		.PKT_CACHE_H               (112),
		.PKT_CACHE_L               (109),
		.PKT_DATA_SIDEBAND_H       (100),
		.PKT_DATA_SIDEBAND_L       (100),
		.PKT_QOS_H                 (102),
		.PKT_QOS_L                 (102),
		.PKT_ADDR_SIDEBAND_H       (99),
		.PKT_ADDR_SIDEBAND_L       (95),
		.PKT_RESPONSE_STATUS_H     (114),
		.PKT_RESPONSE_STATUS_L     (113),
		.ST_DATA_W                 (115),
		.ST_CHANNEL_W              (2),
		.AV_BURSTCOUNT_W           (3),
		.SUPPRESS_0_BYTEEN_RSP     (1),
		.ID                        (0),
		.BURSTWRAP_VALUE           (255),
		.CACHE_VALUE               (0),
		.SECURE_ACCESS_BIT         (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) master_secure_master_translator_avalon_universal_master_0_agent (
		.clk                     (clk_clk),                                                                          //       clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                   // clk_reset.reset
		.av_address              (master_secure_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write                (master_secure_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read                 (master_secure_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata            (master_secure_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata             (master_secure_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest          (master_secure_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid        (master_secure_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable           (master_secure_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount           (master_secure_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess          (master_secure_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock                 (master_secure_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid                (master_secure_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data                 (master_secure_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket        (master_secure_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket          (master_secure_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready                (master_secure_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid                (limiter_rsp_src_valid),                                                            //        rp.valid
		.rp_data                 (limiter_rsp_src_data),                                                             //          .data
		.rp_channel              (limiter_rsp_src_channel),                                                          //          .channel
		.rp_startofpacket        (limiter_rsp_src_startofpacket),                                                    //          .startofpacket
		.rp_endofpacket          (limiter_rsp_src_endofpacket),                                                      //          .endofpacket
		.rp_ready                (limiter_rsp_src_ready),                                                            //          .ready
		.av_response             (),                                                                                 // (terminated)
		.av_writeresponserequest (1'b0),                                                                             // (terminated)
		.av_writeresponsevalid   ()                                                                                  // (terminated)
	);

	altera_merlin_axi_slave_ni #(
		.PKT_QOS_H                   (138),
		.PKT_QOS_L                   (138),
		.PKT_THREAD_ID_H             (141),
		.PKT_THREAD_ID_L             (141),
		.PKT_RESPONSE_STATUS_H       (150),
		.PKT_RESPONSE_STATUS_L       (149),
		.PKT_BEGIN_BURST             (137),
		.PKT_CACHE_H                 (148),
		.PKT_CACHE_L                 (145),
		.PKT_DATA_SIDEBAND_H         (136),
		.PKT_DATA_SIDEBAND_L         (136),
		.PKT_ADDR_SIDEBAND_H         (135),
		.PKT_ADDR_SIDEBAND_L         (131),
		.PKT_BURST_TYPE_H            (130),
		.PKT_BURST_TYPE_L            (129),
		.PKT_PROTECTION_H            (144),
		.PKT_PROTECTION_L            (142),
		.PKT_BURST_SIZE_H            (128),
		.PKT_BURST_SIZE_L            (126),
		.PKT_BURSTWRAP_H             (125),
		.PKT_BURSTWRAP_L             (118),
		.PKT_BYTE_CNT_H              (117),
		.PKT_BYTE_CNT_L              (110),
		.PKT_ADDR_H                  (103),
		.PKT_ADDR_L                  (72),
		.PKT_TRANS_EXCLUSIVE         (109),
		.PKT_TRANS_LOCK              (108),
		.PKT_TRANS_COMPRESSED_READ   (104),
		.PKT_TRANS_POSTED            (105),
		.PKT_TRANS_WRITE             (106),
		.PKT_TRANS_READ              (107),
		.PKT_DATA_H                  (63),
		.PKT_DATA_L                  (0),
		.PKT_BYTEEN_H                (71),
		.PKT_BYTEEN_L                (64),
		.PKT_SRC_ID_H                (139),
		.PKT_SRC_ID_L                (139),
		.PKT_DEST_ID_H               (140),
		.PKT_DEST_ID_L               (140),
		.ADDR_USER_WIDTH             (5),
		.DATA_USER_WIDTH             (1),
		.ST_DATA_W                   (151),
		.ADDR_WIDTH                  (32),
		.RDATA_WIDTH                 (64),
		.WDATA_WIDTH                 (64),
		.ST_CHANNEL_W                (2),
		.AXI_SLAVE_ID_W              (8),
		.PASS_ID_TO_SLAVE            (1),
		.AXI_VERSION                 ("AXI3"),
		.WRITE_ACCEPTANCE_CAPABILITY (8),
		.READ_ACCEPTANCE_CAPABILITY  (8)
	) hps_0_f2h_axi_slave_agent (
		.aclk                   (clk_clk),                                             //        clock_sink.clk
		.aresetn                (~rst_controller_004_reset_out_reset),                 //        reset_sink.reset_n
		.read_cp_valid          (width_adapter_001_cmd_source_valid),                  //           read_cp.valid
		.read_cp_ready          (width_adapter_001_cmd_source_ready),                  //                  .ready
		.read_cp_data           (width_adapter_001_cmd_source_data),                   //                  .data
		.read_cp_channel        (width_adapter_001_cmd_source_channel),                //                  .channel
		.read_cp_startofpacket  (width_adapter_001_cmd_source_startofpacket),          //                  .startofpacket
		.read_cp_endofpacket    (width_adapter_001_cmd_source_endofpacket),            //                  .endofpacket
		.write_cp_ready         (width_adapter_cmd_source_ready),                      //          write_cp.ready
		.write_cp_valid         (width_adapter_cmd_source_valid),                      //                  .valid
		.write_cp_data          (width_adapter_cmd_source_data),                       //                  .data
		.write_cp_channel       (width_adapter_cmd_source_channel),                    //                  .channel
		.write_cp_startofpacket (width_adapter_cmd_source_startofpacket),              //                  .startofpacket
		.write_cp_endofpacket   (width_adapter_cmd_source_endofpacket),                //                  .endofpacket
		.read_rp_ready          (hps_0_f2h_axi_slave_agent_read_rp_ready),             //           read_rp.ready
		.read_rp_valid          (hps_0_f2h_axi_slave_agent_read_rp_valid),             //                  .valid
		.read_rp_data           (hps_0_f2h_axi_slave_agent_read_rp_data),              //                  .data
		.read_rp_startofpacket  (hps_0_f2h_axi_slave_agent_read_rp_startofpacket),     //                  .startofpacket
		.read_rp_endofpacket    (hps_0_f2h_axi_slave_agent_read_rp_endofpacket),       //                  .endofpacket
		.write_rp_ready         (hps_0_f2h_axi_slave_agent_write_rp_ready),            //          write_rp.ready
		.write_rp_valid         (hps_0_f2h_axi_slave_agent_write_rp_valid),            //                  .valid
		.write_rp_data          (hps_0_f2h_axi_slave_agent_write_rp_data),             //                  .data
		.write_rp_startofpacket (hps_0_f2h_axi_slave_agent_write_rp_startofpacket),    //                  .startofpacket
		.write_rp_endofpacket   (hps_0_f2h_axi_slave_agent_write_rp_endofpacket),      //                  .endofpacket
		.awid                   (hps_0_f2h_axi_slave_agent_altera_axi_master_awid),    // altera_axi_master.awid
		.awaddr                 (hps_0_f2h_axi_slave_agent_altera_axi_master_awaddr),  //                  .awaddr
		.awlen                  (hps_0_f2h_axi_slave_agent_altera_axi_master_awlen),   //                  .awlen
		.awsize                 (hps_0_f2h_axi_slave_agent_altera_axi_master_awsize),  //                  .awsize
		.awburst                (hps_0_f2h_axi_slave_agent_altera_axi_master_awburst), //                  .awburst
		.awlock                 (hps_0_f2h_axi_slave_agent_altera_axi_master_awlock),  //                  .awlock
		.awcache                (hps_0_f2h_axi_slave_agent_altera_axi_master_awcache), //                  .awcache
		.awprot                 (hps_0_f2h_axi_slave_agent_altera_axi_master_awprot),  //                  .awprot
		.awuser                 (hps_0_f2h_axi_slave_agent_altera_axi_master_awuser),  //                  .awuser
		.awvalid                (hps_0_f2h_axi_slave_agent_altera_axi_master_awvalid), //                  .awvalid
		.awready                (hps_0_f2h_axi_slave_agent_altera_axi_master_awready), //                  .awready
		.wid                    (hps_0_f2h_axi_slave_agent_altera_axi_master_wid),     //                  .wid
		.wdata                  (hps_0_f2h_axi_slave_agent_altera_axi_master_wdata),   //                  .wdata
		.wstrb                  (hps_0_f2h_axi_slave_agent_altera_axi_master_wstrb),   //                  .wstrb
		.wlast                  (hps_0_f2h_axi_slave_agent_altera_axi_master_wlast),   //                  .wlast
		.wvalid                 (hps_0_f2h_axi_slave_agent_altera_axi_master_wvalid),  //                  .wvalid
		.wready                 (hps_0_f2h_axi_slave_agent_altera_axi_master_wready),  //                  .wready
		.bid                    (hps_0_f2h_axi_slave_agent_altera_axi_master_bid),     //                  .bid
		.bresp                  (hps_0_f2h_axi_slave_agent_altera_axi_master_bresp),   //                  .bresp
		.bvalid                 (hps_0_f2h_axi_slave_agent_altera_axi_master_bvalid),  //                  .bvalid
		.bready                 (hps_0_f2h_axi_slave_agent_altera_axi_master_bready),  //                  .bready
		.arid                   (hps_0_f2h_axi_slave_agent_altera_axi_master_arid),    //                  .arid
		.araddr                 (hps_0_f2h_axi_slave_agent_altera_axi_master_araddr),  //                  .araddr
		.arlen                  (hps_0_f2h_axi_slave_agent_altera_axi_master_arlen),   //                  .arlen
		.arsize                 (hps_0_f2h_axi_slave_agent_altera_axi_master_arsize),  //                  .arsize
		.arburst                (hps_0_f2h_axi_slave_agent_altera_axi_master_arburst), //                  .arburst
		.arlock                 (hps_0_f2h_axi_slave_agent_altera_axi_master_arlock),  //                  .arlock
		.arcache                (hps_0_f2h_axi_slave_agent_altera_axi_master_arcache), //                  .arcache
		.arprot                 (hps_0_f2h_axi_slave_agent_altera_axi_master_arprot),  //                  .arprot
		.aruser                 (hps_0_f2h_axi_slave_agent_altera_axi_master_aruser),  //                  .aruser
		.arvalid                (hps_0_f2h_axi_slave_agent_altera_axi_master_arvalid), //                  .arvalid
		.arready                (hps_0_f2h_axi_slave_agent_altera_axi_master_arready), //                  .arready
		.rid                    (hps_0_f2h_axi_slave_agent_altera_axi_master_rid),     //                  .rid
		.rdata                  (hps_0_f2h_axi_slave_agent_altera_axi_master_rdata),   //                  .rdata
		.rresp                  (hps_0_f2h_axi_slave_agent_altera_axi_master_rresp),   //                  .rresp
		.rlast                  (hps_0_f2h_axi_slave_agent_altera_axi_master_rlast),   //                  .rlast
		.rvalid                 (hps_0_f2h_axi_slave_agent_altera_axi_master_rvalid),  //                  .rvalid
		.rready                 (hps_0_f2h_axi_slave_agent_altera_axi_master_rready)   //                  .rready
	);

	altera_merlin_axi_master_ni #(
		.ID_WIDTH                  (12),
		.ADDR_WIDTH                (21),
		.RDATA_WIDTH               (32),
		.WDATA_WIDTH               (32),
		.ADDR_USER_WIDTH           (1),
		.DATA_USER_WIDTH           (1),
		.AXI_BURST_LENGTH_WIDTH    (4),
		.AXI_LOCK_WIDTH            (2),
		.AXI_VERSION               ("AXI3"),
		.WRITE_ISSUING_CAPABILITY  (8),
		.READ_ISSUING_CAPABILITY   (8),
		.PKT_BEGIN_BURST           (84),
		.PKT_CACHE_H               (110),
		.PKT_CACHE_L               (107),
		.PKT_ADDR_SIDEBAND_H       (82),
		.PKT_ADDR_SIDEBAND_L       (82),
		.PKT_PROTECTION_H          (106),
		.PKT_PROTECTION_L          (104),
		.PKT_BURST_SIZE_H          (79),
		.PKT_BURST_SIZE_L          (77),
		.PKT_BURST_TYPE_H          (81),
		.PKT_BURST_TYPE_L          (80),
		.PKT_RESPONSE_STATUS_L     (111),
		.PKT_RESPONSE_STATUS_H     (112),
		.PKT_BURSTWRAP_H           (76),
		.PKT_BURSTWRAP_L           (70),
		.PKT_BYTE_CNT_H            (69),
		.PKT_BYTE_CNT_L            (63),
		.PKT_ADDR_H                (56),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_EXCLUSIVE       (62),
		.PKT_TRANS_LOCK            (61),
		.PKT_TRANS_COMPRESSED_READ (57),
		.PKT_TRANS_POSTED          (58),
		.PKT_TRANS_WRITE           (59),
		.PKT_TRANS_READ            (60),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (88),
		.PKT_SRC_ID_L              (86),
		.PKT_DEST_ID_H             (91),
		.PKT_DEST_ID_L             (89),
		.PKT_THREAD_ID_H           (103),
		.PKT_THREAD_ID_L           (92),
		.PKT_QOS_L                 (85),
		.PKT_QOS_H                 (85),
		.PKT_DATA_SIDEBAND_H       (83),
		.PKT_DATA_SIDEBAND_L       (83),
		.ST_DATA_W                 (113),
		.ST_CHANNEL_W              (8),
		.ID                        (0)
	) hps_0_h2f_lw_axi_master_agent (
		.aclk                   (clk_clk),                                              //              clk.clk
		.aresetn                (~rst_controller_004_reset_out_reset),                  //        clk_reset.reset_n
		.write_cp_valid         (hps_0_h2f_lw_axi_master_agent_write_cp_valid),         //         write_cp.valid
		.write_cp_data          (hps_0_h2f_lw_axi_master_agent_write_cp_data),          //                 .data
		.write_cp_startofpacket (hps_0_h2f_lw_axi_master_agent_write_cp_startofpacket), //                 .startofpacket
		.write_cp_endofpacket   (hps_0_h2f_lw_axi_master_agent_write_cp_endofpacket),   //                 .endofpacket
		.write_cp_ready         (hps_0_h2f_lw_axi_master_agent_write_cp_ready),         //                 .ready
		.write_rp_valid         (limiter_001_rsp_src_valid),                            //         write_rp.valid
		.write_rp_data          (limiter_001_rsp_src_data),                             //                 .data
		.write_rp_channel       (limiter_001_rsp_src_channel),                          //                 .channel
		.write_rp_startofpacket (limiter_001_rsp_src_startofpacket),                    //                 .startofpacket
		.write_rp_endofpacket   (limiter_001_rsp_src_endofpacket),                      //                 .endofpacket
		.write_rp_ready         (limiter_001_rsp_src_ready),                            //                 .ready
		.read_cp_valid          (hps_0_h2f_lw_axi_master_agent_read_cp_valid),          //          read_cp.valid
		.read_cp_data           (hps_0_h2f_lw_axi_master_agent_read_cp_data),           //                 .data
		.read_cp_startofpacket  (hps_0_h2f_lw_axi_master_agent_read_cp_startofpacket),  //                 .startofpacket
		.read_cp_endofpacket    (hps_0_h2f_lw_axi_master_agent_read_cp_endofpacket),    //                 .endofpacket
		.read_cp_ready          (hps_0_h2f_lw_axi_master_agent_read_cp_ready),          //                 .ready
		.read_rp_valid          (limiter_002_rsp_src_valid),                            //          read_rp.valid
		.read_rp_data           (limiter_002_rsp_src_data),                             //                 .data
		.read_rp_channel        (limiter_002_rsp_src_channel),                          //                 .channel
		.read_rp_startofpacket  (limiter_002_rsp_src_startofpacket),                    //                 .startofpacket
		.read_rp_endofpacket    (limiter_002_rsp_src_endofpacket),                      //                 .endofpacket
		.read_rp_ready          (limiter_002_rsp_src_ready),                            //                 .ready
		.awid                   (hps_0_h2f_lw_axi_master_awid),                         // altera_axi_slave.awid
		.awaddr                 (hps_0_h2f_lw_axi_master_awaddr),                       //                 .awaddr
		.awlen                  (hps_0_h2f_lw_axi_master_awlen),                        //                 .awlen
		.awsize                 (hps_0_h2f_lw_axi_master_awsize),                       //                 .awsize
		.awburst                (hps_0_h2f_lw_axi_master_awburst),                      //                 .awburst
		.awlock                 (hps_0_h2f_lw_axi_master_awlock),                       //                 .awlock
		.awcache                (hps_0_h2f_lw_axi_master_awcache),                      //                 .awcache
		.awprot                 (hps_0_h2f_lw_axi_master_awprot),                       //                 .awprot
		.awvalid                (hps_0_h2f_lw_axi_master_awvalid),                      //                 .awvalid
		.awready                (hps_0_h2f_lw_axi_master_awready),                      //                 .awready
		.wid                    (hps_0_h2f_lw_axi_master_wid),                          //                 .wid
		.wdata                  (hps_0_h2f_lw_axi_master_wdata),                        //                 .wdata
		.wstrb                  (hps_0_h2f_lw_axi_master_wstrb),                        //                 .wstrb
		.wlast                  (hps_0_h2f_lw_axi_master_wlast),                        //                 .wlast
		.wvalid                 (hps_0_h2f_lw_axi_master_wvalid),                       //                 .wvalid
		.wready                 (hps_0_h2f_lw_axi_master_wready),                       //                 .wready
		.bid                    (hps_0_h2f_lw_axi_master_bid),                          //                 .bid
		.bresp                  (hps_0_h2f_lw_axi_master_bresp),                        //                 .bresp
		.bvalid                 (hps_0_h2f_lw_axi_master_bvalid),                       //                 .bvalid
		.bready                 (hps_0_h2f_lw_axi_master_bready),                       //                 .bready
		.arid                   (hps_0_h2f_lw_axi_master_arid),                         //                 .arid
		.araddr                 (hps_0_h2f_lw_axi_master_araddr),                       //                 .araddr
		.arlen                  (hps_0_h2f_lw_axi_master_arlen),                        //                 .arlen
		.arsize                 (hps_0_h2f_lw_axi_master_arsize),                       //                 .arsize
		.arburst                (hps_0_h2f_lw_axi_master_arburst),                      //                 .arburst
		.arlock                 (hps_0_h2f_lw_axi_master_arlock),                       //                 .arlock
		.arcache                (hps_0_h2f_lw_axi_master_arcache),                      //                 .arcache
		.arprot                 (hps_0_h2f_lw_axi_master_arprot),                       //                 .arprot
		.arvalid                (hps_0_h2f_lw_axi_master_arvalid),                      //                 .arvalid
		.arready                (hps_0_h2f_lw_axi_master_arready),                      //                 .arready
		.rid                    (hps_0_h2f_lw_axi_master_rid),                          //                 .rid
		.rdata                  (hps_0_h2f_lw_axi_master_rdata),                        //                 .rdata
		.rresp                  (hps_0_h2f_lw_axi_master_rresp),                        //                 .rresp
		.rlast                  (hps_0_h2f_lw_axi_master_rlast),                        //                 .rlast
		.rvalid                 (hps_0_h2f_lw_axi_master_rvalid),                       //                 .rvalid
		.rready                 (hps_0_h2f_lw_axi_master_rready),                       //                 .rready
		.awuser                 (1'b0),                                                 //      (terminated)
		.aruser                 (1'b0),                                                 //      (terminated)
		.awqos                  (4'b0000),                                              //      (terminated)
		.arqos                  (4'b0000),                                              //      (terminated)
		.awregion               (4'b0000),                                              //      (terminated)
		.arregion               (4'b0000),                                              //      (terminated)
		.wuser                  (1'b0),                                                 //      (terminated)
		.ruser                  (),                                                     //      (terminated)
		.buser                  ()                                                      //      (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (84),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (56),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (57),
		.PKT_TRANS_POSTED          (58),
		.PKT_TRANS_WRITE           (59),
		.PKT_TRANS_READ            (60),
		.PKT_TRANS_LOCK            (61),
		.PKT_SRC_ID_H              (88),
		.PKT_SRC_ID_L              (86),
		.PKT_DEST_ID_H             (91),
		.PKT_DEST_ID_L             (89),
		.PKT_BURSTWRAP_H           (76),
		.PKT_BURSTWRAP_L           (70),
		.PKT_BYTE_CNT_H            (69),
		.PKT_BYTE_CNT_L            (63),
		.PKT_PROTECTION_H          (106),
		.PKT_PROTECTION_L          (104),
		.PKT_RESPONSE_STATUS_H     (112),
		.PKT_RESPONSE_STATUS_L     (111),
		.PKT_BURST_SIZE_H          (79),
		.PKT_BURST_SIZE_L          (77),
		.ST_CHANNEL_W              (8),
		.ST_DATA_W                 (113),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) led_pio_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                         //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                  //       clk_reset.reset
		.m0_address              (led_pio_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (led_pio_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (led_pio_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (led_pio_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (led_pio_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (led_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (led_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (led_pio_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (led_pio_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (led_pio_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (led_pio_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (led_pio_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (led_pio_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (led_pio_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (led_pio_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (led_pio_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_source0_ready),                                                     //              cp.ready
		.cp_valid                (burst_adapter_source0_valid),                                                     //                .valid
		.cp_data                 (burst_adapter_source0_data),                                                      //                .data
		.cp_startofpacket        (burst_adapter_source0_startofpacket),                                             //                .startofpacket
		.cp_endofpacket          (burst_adapter_source0_endofpacket),                                               //                .endofpacket
		.cp_channel              (burst_adapter_source0_channel),                                                   //                .channel
		.rf_sink_ready           (led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (led_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (led_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (led_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (led_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (led_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                           //     (terminated)
		.m0_writeresponserequest (),                                                                                //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                             //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (114),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                         //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                  // clk_reset.reset
		.in_data           (led_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (led_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (led_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (led_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (led_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (led_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                           // (terminated)
		.csr_read          (1'b0),                                                                            // (terminated)
		.csr_write         (1'b0),                                                                            // (terminated)
		.csr_readdata      (),                                                                                // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                            // (terminated)
		.almost_full_data  (),                                                                                // (terminated)
		.almost_empty_data (),                                                                                // (terminated)
		.in_empty          (1'b0),                                                                            // (terminated)
		.out_empty         (),                                                                                // (terminated)
		.in_error          (1'b0),                                                                            // (terminated)
		.out_error         (),                                                                                // (terminated)
		.in_channel        (1'b0),                                                                            // (terminated)
		.out_channel       ()                                                                                 // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (34),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (clk_clk),                                                                   //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                            // clk_reset.reset
		.in_data           (led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (led_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                     // (terminated)
		.csr_read          (1'b0),                                                                      // (terminated)
		.csr_write         (1'b0),                                                                      // (terminated)
		.csr_readdata      (),                                                                          // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                      // (terminated)
		.almost_full_data  (),                                                                          // (terminated)
		.almost_empty_data (),                                                                          // (terminated)
		.in_startofpacket  (1'b0),                                                                      // (terminated)
		.in_endofpacket    (1'b0),                                                                      // (terminated)
		.out_startofpacket (),                                                                          // (terminated)
		.out_endofpacket   (),                                                                          // (terminated)
		.in_empty          (1'b0),                                                                      // (terminated)
		.out_empty         (),                                                                          // (terminated)
		.in_error          (1'b0),                                                                      // (terminated)
		.out_error         (),                                                                          // (terminated)
		.in_channel        (1'b0),                                                                      // (terminated)
		.out_channel       ()                                                                           // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (84),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (56),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (57),
		.PKT_TRANS_POSTED          (58),
		.PKT_TRANS_WRITE           (59),
		.PKT_TRANS_READ            (60),
		.PKT_TRANS_LOCK            (61),
		.PKT_SRC_ID_H              (88),
		.PKT_SRC_ID_L              (86),
		.PKT_DEST_ID_H             (91),
		.PKT_DEST_ID_L             (89),
		.PKT_BURSTWRAP_H           (76),
		.PKT_BURSTWRAP_L           (70),
		.PKT_BYTE_CNT_H            (69),
		.PKT_BYTE_CNT_L            (63),
		.PKT_PROTECTION_H          (106),
		.PKT_PROTECTION_L          (104),
		.PKT_RESPONSE_STATUS_H     (112),
		.PKT_RESPONSE_STATUS_L     (111),
		.PKT_BURST_SIZE_H          (79),
		.PKT_BURST_SIZE_L          (77),
		.ST_CHANNEL_W              (8),
		.ST_DATA_W                 (113),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) dipsw_pio_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                           //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                    //       clk_reset.reset
		.m0_address              (dipsw_pio_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (dipsw_pio_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (dipsw_pio_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (dipsw_pio_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (dipsw_pio_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (dipsw_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (dipsw_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (dipsw_pio_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (dipsw_pio_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (dipsw_pio_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (dipsw_pio_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (dipsw_pio_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (dipsw_pio_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (dipsw_pio_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (dipsw_pio_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (dipsw_pio_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_001_source0_ready),                                                   //              cp.ready
		.cp_valid                (burst_adapter_001_source0_valid),                                                   //                .valid
		.cp_data                 (burst_adapter_001_source0_data),                                                    //                .data
		.cp_startofpacket        (burst_adapter_001_source0_startofpacket),                                           //                .startofpacket
		.cp_endofpacket          (burst_adapter_001_source0_endofpacket),                                             //                .endofpacket
		.cp_channel              (burst_adapter_001_source0_channel),                                                 //                .channel
		.rf_sink_ready           (dipsw_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (dipsw_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (dipsw_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (dipsw_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (dipsw_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (dipsw_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (dipsw_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (dipsw_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (dipsw_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (dipsw_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (dipsw_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (dipsw_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (dipsw_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (dipsw_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (dipsw_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (dipsw_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                             //     (terminated)
		.m0_writeresponserequest (),                                                                                  //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                               //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (114),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) dipsw_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                           //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                    // clk_reset.reset
		.in_data           (dipsw_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (dipsw_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (dipsw_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (dipsw_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (dipsw_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (dipsw_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (dipsw_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (dipsw_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (dipsw_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (dipsw_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                             // (terminated)
		.csr_read          (1'b0),                                                                              // (terminated)
		.csr_write         (1'b0),                                                                              // (terminated)
		.csr_readdata      (),                                                                                  // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                              // (terminated)
		.almost_full_data  (),                                                                                  // (terminated)
		.almost_empty_data (),                                                                                  // (terminated)
		.in_empty          (1'b0),                                                                              // (terminated)
		.out_empty         (),                                                                                  // (terminated)
		.in_error          (1'b0),                                                                              // (terminated)
		.out_error         (),                                                                                  // (terminated)
		.in_channel        (1'b0),                                                                              // (terminated)
		.out_channel       ()                                                                                   // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (34),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) dipsw_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (clk_clk),                                                                     //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                              // clk_reset.reset
		.in_data           (dipsw_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (dipsw_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (dipsw_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (dipsw_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (dipsw_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (dipsw_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                       // (terminated)
		.csr_read          (1'b0),                                                                        // (terminated)
		.csr_write         (1'b0),                                                                        // (terminated)
		.csr_readdata      (),                                                                            // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                        // (terminated)
		.almost_full_data  (),                                                                            // (terminated)
		.almost_empty_data (),                                                                            // (terminated)
		.in_startofpacket  (1'b0),                                                                        // (terminated)
		.in_endofpacket    (1'b0),                                                                        // (terminated)
		.out_startofpacket (),                                                                            // (terminated)
		.out_endofpacket   (),                                                                            // (terminated)
		.in_empty          (1'b0),                                                                        // (terminated)
		.out_empty         (),                                                                            // (terminated)
		.in_error          (1'b0),                                                                        // (terminated)
		.out_error         (),                                                                            // (terminated)
		.in_channel        (1'b0),                                                                        // (terminated)
		.out_channel       ()                                                                             // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (84),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (56),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (57),
		.PKT_TRANS_POSTED          (58),
		.PKT_TRANS_WRITE           (59),
		.PKT_TRANS_READ            (60),
		.PKT_TRANS_LOCK            (61),
		.PKT_SRC_ID_H              (88),
		.PKT_SRC_ID_L              (86),
		.PKT_DEST_ID_H             (91),
		.PKT_DEST_ID_L             (89),
		.PKT_BURSTWRAP_H           (76),
		.PKT_BURSTWRAP_L           (70),
		.PKT_BYTE_CNT_H            (69),
		.PKT_BYTE_CNT_L            (63),
		.PKT_PROTECTION_H          (106),
		.PKT_PROTECTION_L          (104),
		.PKT_RESPONSE_STATUS_H     (112),
		.PKT_RESPONSE_STATUS_L     (111),
		.PKT_BURST_SIZE_H          (79),
		.PKT_BURST_SIZE_L          (77),
		.ST_CHANNEL_W              (8),
		.ST_DATA_W                 (113),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) button_pio_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                            //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                     //       clk_reset.reset
		.m0_address              (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (button_pio_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (button_pio_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (button_pio_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (button_pio_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (button_pio_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (button_pio_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_002_source0_ready),                                                    //              cp.ready
		.cp_valid                (burst_adapter_002_source0_valid),                                                    //                .valid
		.cp_data                 (burst_adapter_002_source0_data),                                                     //                .data
		.cp_startofpacket        (burst_adapter_002_source0_startofpacket),                                            //                .startofpacket
		.cp_endofpacket          (burst_adapter_002_source0_endofpacket),                                              //                .endofpacket
		.cp_channel              (burst_adapter_002_source0_channel),                                                  //                .channel
		.rf_sink_ready           (button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (button_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (button_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (button_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (button_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (button_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (button_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (button_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (button_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (button_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (button_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (button_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                              //     (terminated)
		.m0_writeresponserequest (),                                                                                   //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (114),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                            //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                     // clk_reset.reset
		.in_data           (button_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (button_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (button_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (button_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (button_pio_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (button_pio_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                              // (terminated)
		.csr_read          (1'b0),                                                                               // (terminated)
		.csr_write         (1'b0),                                                                               // (terminated)
		.csr_readdata      (),                                                                                   // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                               // (terminated)
		.almost_full_data  (),                                                                                   // (terminated)
		.almost_empty_data (),                                                                                   // (terminated)
		.in_empty          (1'b0),                                                                               // (terminated)
		.out_empty         (),                                                                                   // (terminated)
		.in_error          (1'b0),                                                                               // (terminated)
		.out_error         (),                                                                                   // (terminated)
		.in_channel        (1'b0),                                                                               // (terminated)
		.out_channel       ()                                                                                    // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (34),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) button_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (clk_clk),                                                                      //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                               // clk_reset.reset
		.in_data           (button_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (button_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (button_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (button_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (button_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (button_pio_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                        // (terminated)
		.csr_read          (1'b0),                                                                         // (terminated)
		.csr_write         (1'b0),                                                                         // (terminated)
		.csr_readdata      (),                                                                             // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                         // (terminated)
		.almost_full_data  (),                                                                             // (terminated)
		.almost_empty_data (),                                                                             // (terminated)
		.in_startofpacket  (1'b0),                                                                         // (terminated)
		.in_endofpacket    (1'b0),                                                                         // (terminated)
		.out_startofpacket (),                                                                             // (terminated)
		.out_endofpacket   (),                                                                             // (terminated)
		.in_empty          (1'b0),                                                                         // (terminated)
		.out_empty         (),                                                                             // (terminated)
		.in_error          (1'b0),                                                                         // (terminated)
		.out_error         (),                                                                             // (terminated)
		.in_channel        (1'b0),                                                                         // (terminated)
		.out_channel       ()                                                                              // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (84),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (56),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (57),
		.PKT_TRANS_POSTED          (58),
		.PKT_TRANS_WRITE           (59),
		.PKT_TRANS_READ            (60),
		.PKT_TRANS_LOCK            (61),
		.PKT_SRC_ID_H              (88),
		.PKT_SRC_ID_L              (86),
		.PKT_DEST_ID_H             (91),
		.PKT_DEST_ID_L             (89),
		.PKT_BURSTWRAP_H           (76),
		.PKT_BURSTWRAP_L           (70),
		.PKT_BYTE_CNT_H            (69),
		.PKT_BYTE_CNT_L            (63),
		.PKT_PROTECTION_H          (106),
		.PKT_PROTECTION_L          (104),
		.PKT_RESPONSE_STATUS_H     (112),
		.PKT_RESPONSE_STATUS_L     (111),
		.PKT_BURST_SIZE_H          (79),
		.PKT_BURST_SIZE_L          (77),
		.ST_CHANNEL_W              (8),
		.ST_DATA_W                 (113),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                          //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                   //       clk_reset.reset
		.m0_address              (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_003_source0_ready),                                                                  //              cp.ready
		.cp_valid                (burst_adapter_003_source0_valid),                                                                  //                .valid
		.cp_data                 (burst_adapter_003_source0_data),                                                                   //                .data
		.cp_startofpacket        (burst_adapter_003_source0_startofpacket),                                                          //                .startofpacket
		.cp_endofpacket          (burst_adapter_003_source0_endofpacket),                                                            //                .endofpacket
		.cp_channel              (burst_adapter_003_source0_channel),                                                                //                .channel
		.rf_sink_ready           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                            //     (terminated)
		.m0_writeresponserequest (),                                                                                                 //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                              //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (114),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                          //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                   // clk_reset.reset
		.in_data           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                            // (terminated)
		.csr_read          (1'b0),                                                                                             // (terminated)
		.csr_write         (1'b0),                                                                                             // (terminated)
		.csr_readdata      (),                                                                                                 // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                             // (terminated)
		.almost_full_data  (),                                                                                                 // (terminated)
		.almost_empty_data (),                                                                                                 // (terminated)
		.in_empty          (1'b0),                                                                                             // (terminated)
		.out_empty         (),                                                                                                 // (terminated)
		.in_error          (1'b0),                                                                                             // (terminated)
		.out_error         (),                                                                                                 // (terminated)
		.in_channel        (1'b0),                                                                                             // (terminated)
		.out_channel       ()                                                                                                  // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (34),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (clk_clk),                                                                                    //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                             // clk_reset.reset
		.in_data           (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                                      // (terminated)
		.csr_read          (1'b0),                                                                                       // (terminated)
		.csr_write         (1'b0),                                                                                       // (terminated)
		.csr_readdata      (),                                                                                           // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                       // (terminated)
		.almost_full_data  (),                                                                                           // (terminated)
		.almost_empty_data (),                                                                                           // (terminated)
		.in_startofpacket  (1'b0),                                                                                       // (terminated)
		.in_endofpacket    (1'b0),                                                                                       // (terminated)
		.out_startofpacket (),                                                                                           // (terminated)
		.out_endofpacket   (),                                                                                           // (terminated)
		.in_empty          (1'b0),                                                                                       // (terminated)
		.out_empty         (),                                                                                           // (terminated)
		.in_error          (1'b0),                                                                                       // (terminated)
		.out_error         (),                                                                                           // (terminated)
		.in_channel        (1'b0),                                                                                       // (terminated)
		.out_channel       ()                                                                                            // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (84),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (56),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (57),
		.PKT_TRANS_POSTED          (58),
		.PKT_TRANS_WRITE           (59),
		.PKT_TRANS_READ            (60),
		.PKT_TRANS_LOCK            (61),
		.PKT_SRC_ID_H              (88),
		.PKT_SRC_ID_L              (86),
		.PKT_DEST_ID_H             (91),
		.PKT_DEST_ID_L             (89),
		.PKT_BURSTWRAP_H           (76),
		.PKT_BURSTWRAP_L           (70),
		.PKT_BYTE_CNT_H            (69),
		.PKT_BYTE_CNT_L            (63),
		.PKT_PROTECTION_H          (106),
		.PKT_PROTECTION_L          (104),
		.PKT_RESPONSE_STATUS_H     (112),
		.PKT_RESPONSE_STATUS_L     (111),
		.PKT_BURST_SIZE_H          (79),
		.PKT_BURST_SIZE_L          (77),
		.ST_CHANNEL_W              (8),
		.ST_DATA_W                 (113),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent (
		.clk                     (clk_clk),                                                                                             //             clk.clk
		.reset                   (rst_controller_reset_out_reset),                                                                      //       clk_reset.reset
		.m0_address              (oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_004_source0_ready),                                                                     //              cp.ready
		.cp_valid                (burst_adapter_004_source0_valid),                                                                     //                .valid
		.cp_data                 (burst_adapter_004_source0_data),                                                                      //                .data
		.cp_startofpacket        (burst_adapter_004_source0_startofpacket),                                                             //                .startofpacket
		.cp_endofpacket          (burst_adapter_004_source0_endofpacket),                                                               //                .endofpacket
		.cp_channel              (burst_adapter_004_source0_channel),                                                                   //                .channel
		.rf_sink_ready           (oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                               //     (terminated)
		.m0_writeresponserequest (),                                                                                                    //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                                 //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (114),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (clk_clk),                                                                                             //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                      // clk_reset.reset
		.in_data           (oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                               // (terminated)
		.csr_read          (1'b0),                                                                                                // (terminated)
		.csr_write         (1'b0),                                                                                                // (terminated)
		.csr_readdata      (),                                                                                                    // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                                // (terminated)
		.almost_full_data  (),                                                                                                    // (terminated)
		.almost_empty_data (),                                                                                                    // (terminated)
		.in_empty          (1'b0),                                                                                                // (terminated)
		.out_empty         (),                                                                                                    // (terminated)
		.in_error          (1'b0),                                                                                                // (terminated)
		.out_error         (),                                                                                                    // (terminated)
		.in_channel        (1'b0),                                                                                                // (terminated)
		.out_channel       ()                                                                                                     // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (34),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (clk_clk),                                                                                       //       clk.clk
		.reset             (rst_controller_reset_out_reset),                                                                // clk_reset.reset
		.in_data           (oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                                         // (terminated)
		.csr_read          (1'b0),                                                                                          // (terminated)
		.csr_write         (1'b0),                                                                                          // (terminated)
		.csr_readdata      (),                                                                                              // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                          // (terminated)
		.almost_full_data  (),                                                                                              // (terminated)
		.almost_empty_data (),                                                                                              // (terminated)
		.in_startofpacket  (1'b0),                                                                                          // (terminated)
		.in_endofpacket    (1'b0),                                                                                          // (terminated)
		.out_startofpacket (),                                                                                              // (terminated)
		.out_endofpacket   (),                                                                                              // (terminated)
		.in_empty          (1'b0),                                                                                          // (terminated)
		.out_empty         (),                                                                                              // (terminated)
		.in_error          (1'b0),                                                                                          // (terminated)
		.out_error         (),                                                                                              // (terminated)
		.in_channel        (1'b0),                                                                                          // (terminated)
		.out_channel       ()                                                                                               // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (84),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (56),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (57),
		.PKT_TRANS_POSTED          (58),
		.PKT_TRANS_WRITE           (59),
		.PKT_TRANS_READ            (60),
		.PKT_TRANS_LOCK            (61),
		.PKT_SRC_ID_H              (88),
		.PKT_SRC_ID_L              (86),
		.PKT_DEST_ID_H             (91),
		.PKT_DEST_ID_L             (89),
		.PKT_BURSTWRAP_H           (76),
		.PKT_BURSTWRAP_L           (70),
		.PKT_BYTE_CNT_H            (69),
		.PKT_BYTE_CNT_L            (63),
		.PKT_PROTECTION_H          (106),
		.PKT_PROTECTION_L          (104),
		.PKT_RESPONSE_STATUS_H     (112),
		.PKT_RESPONSE_STATUS_L     (111),
		.PKT_BURST_SIZE_H          (79),
		.PKT_BURST_SIZE_L          (77),
		.ST_CHANNEL_W              (8),
		.ST_DATA_W                 (113),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent (
		.clk                     (pll_stream_outclk1_clk),                                                                     //             clk.clk
		.reset                   (rst_controller_002_reset_out_reset),                                                         //       clk_reset.reset
		.m0_address              (alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_005_source0_ready),                                                            //              cp.ready
		.cp_valid                (burst_adapter_005_source0_valid),                                                            //                .valid
		.cp_data                 (burst_adapter_005_source0_data),                                                             //                .data
		.cp_startofpacket        (burst_adapter_005_source0_startofpacket),                                                    //                .startofpacket
		.cp_endofpacket          (burst_adapter_005_source0_endofpacket),                                                      //                .endofpacket
		.cp_channel              (burst_adapter_005_source0_channel),                                                          //                .channel
		.rf_sink_ready           (alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                      //     (terminated)
		.m0_writeresponserequest (),                                                                                           //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                        //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (114),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (pll_stream_outclk1_clk),                                                                     //       clk.clk
		.reset             (rst_controller_002_reset_out_reset),                                                         // clk_reset.reset
		.in_data           (alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                      // (terminated)
		.csr_read          (1'b0),                                                                                       // (terminated)
		.csr_write         (1'b0),                                                                                       // (terminated)
		.csr_readdata      (),                                                                                           // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                       // (terminated)
		.almost_full_data  (),                                                                                           // (terminated)
		.almost_empty_data (),                                                                                           // (terminated)
		.in_empty          (1'b0),                                                                                       // (terminated)
		.out_empty         (),                                                                                           // (terminated)
		.in_error          (1'b0),                                                                                       // (terminated)
		.out_error         (),                                                                                           // (terminated)
		.in_channel        (1'b0),                                                                                       // (terminated)
		.out_channel       ()                                                                                            // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (34),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (pll_stream_outclk1_clk),                                                               //       clk.clk
		.reset             (rst_controller_002_reset_out_reset),                                                   // clk_reset.reset
		.in_data           (alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                                // (terminated)
		.csr_read          (1'b0),                                                                                 // (terminated)
		.csr_write         (1'b0),                                                                                 // (terminated)
		.csr_readdata      (),                                                                                     // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                 // (terminated)
		.almost_full_data  (),                                                                                     // (terminated)
		.almost_empty_data (),                                                                                     // (terminated)
		.in_startofpacket  (1'b0),                                                                                 // (terminated)
		.in_endofpacket    (1'b0),                                                                                 // (terminated)
		.out_startofpacket (),                                                                                     // (terminated)
		.out_endofpacket   (),                                                                                     // (terminated)
		.in_empty          (1'b0),                                                                                 // (terminated)
		.out_empty         (),                                                                                     // (terminated)
		.in_error          (1'b0),                                                                                 // (terminated)
		.out_error         (),                                                                                     // (terminated)
		.in_channel        (1'b0),                                                                                 // (terminated)
		.out_channel       ()                                                                                      // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (84),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (56),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (57),
		.PKT_TRANS_POSTED          (58),
		.PKT_TRANS_WRITE           (59),
		.PKT_TRANS_READ            (60),
		.PKT_TRANS_LOCK            (61),
		.PKT_SRC_ID_H              (88),
		.PKT_SRC_ID_L              (86),
		.PKT_DEST_ID_H             (91),
		.PKT_DEST_ID_L             (89),
		.PKT_BURSTWRAP_H           (76),
		.PKT_BURSTWRAP_L           (70),
		.PKT_BYTE_CNT_H            (69),
		.PKT_BYTE_CNT_L            (63),
		.PKT_PROTECTION_H          (106),
		.PKT_PROTECTION_L          (104),
		.PKT_RESPONSE_STATUS_H     (112),
		.PKT_RESPONSE_STATUS_L     (111),
		.PKT_BURST_SIZE_H          (79),
		.PKT_BURST_SIZE_L          (77),
		.ST_CHANNEL_W              (8),
		.ST_DATA_W                 (113),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (pll_stream_outclk1_clk),                                                                          //             clk.clk
		.reset                   (rst_controller_002_reset_out_reset),                                                              //       clk_reset.reset
		.m0_address              (alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_006_source0_ready),                                                                 //              cp.ready
		.cp_valid                (burst_adapter_006_source0_valid),                                                                 //                .valid
		.cp_data                 (burst_adapter_006_source0_data),                                                                  //                .data
		.cp_startofpacket        (burst_adapter_006_source0_startofpacket),                                                         //                .startofpacket
		.cp_endofpacket          (burst_adapter_006_source0_endofpacket),                                                           //                .endofpacket
		.cp_channel              (burst_adapter_006_source0_channel),                                                               //                .channel
		.rf_sink_ready           (alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                           //     (terminated)
		.m0_writeresponserequest (),                                                                                                //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                             //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (114),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (pll_stream_outclk1_clk),                                                                          //       clk.clk
		.reset             (rst_controller_002_reset_out_reset),                                                              // clk_reset.reset
		.in_data           (alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                           // (terminated)
		.csr_read          (1'b0),                                                                                            // (terminated)
		.csr_write         (1'b0),                                                                                            // (terminated)
		.csr_readdata      (),                                                                                                // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                            // (terminated)
		.almost_full_data  (),                                                                                                // (terminated)
		.almost_empty_data (),                                                                                                // (terminated)
		.in_empty          (1'b0),                                                                                            // (terminated)
		.out_empty         (),                                                                                                // (terminated)
		.in_error          (1'b0),                                                                                            // (terminated)
		.out_error         (),                                                                                                // (terminated)
		.in_channel        (1'b0),                                                                                            // (terminated)
		.out_channel       ()                                                                                                 // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (34),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (pll_stream_outclk1_clk),                                                                    //       clk.clk
		.reset             (rst_controller_002_reset_out_reset),                                                        // clk_reset.reset
		.in_data           (alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                                     // (terminated)
		.csr_read          (1'b0),                                                                                      // (terminated)
		.csr_write         (1'b0),                                                                                      // (terminated)
		.csr_readdata      (),                                                                                          // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                      // (terminated)
		.almost_full_data  (),                                                                                          // (terminated)
		.almost_empty_data (),                                                                                          // (terminated)
		.in_startofpacket  (1'b0),                                                                                      // (terminated)
		.in_endofpacket    (1'b0),                                                                                      // (terminated)
		.out_startofpacket (),                                                                                          // (terminated)
		.out_endofpacket   (),                                                                                          // (terminated)
		.in_empty          (1'b0),                                                                                      // (terminated)
		.out_empty         (),                                                                                          // (terminated)
		.in_error          (1'b0),                                                                                      // (terminated)
		.out_error         (),                                                                                          // (terminated)
		.in_channel        (1'b0),                                                                                      // (terminated)
		.out_channel       ()                                                                                           // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (84),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_ADDR_H                (56),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (57),
		.PKT_TRANS_POSTED          (58),
		.PKT_TRANS_WRITE           (59),
		.PKT_TRANS_READ            (60),
		.PKT_TRANS_LOCK            (61),
		.PKT_SRC_ID_H              (88),
		.PKT_SRC_ID_L              (86),
		.PKT_DEST_ID_H             (91),
		.PKT_DEST_ID_L             (89),
		.PKT_BURSTWRAP_H           (76),
		.PKT_BURSTWRAP_L           (70),
		.PKT_BYTE_CNT_H            (69),
		.PKT_BYTE_CNT_L            (63),
		.PKT_PROTECTION_H          (106),
		.PKT_PROTECTION_L          (104),
		.PKT_RESPONSE_STATUS_H     (112),
		.PKT_RESPONSE_STATUS_L     (111),
		.PKT_BURST_SIZE_H          (79),
		.PKT_BURST_SIZE_L          (77),
		.ST_CHANNEL_W              (8),
		.ST_DATA_W                 (113),
		.AVS_BURSTCOUNT_W          (3),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) audio_if_0_avalon_slave_translator_avalon_universal_slave_0_agent (
		.clk                     (pll_audio_outclk0_clk),                                                                        //             clk.clk
		.reset                   (rst_controller_003_reset_out_reset),                                                           //       clk_reset.reset
		.m0_address              (audio_if_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (audio_if_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (audio_if_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (audio_if_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (audio_if_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (audio_if_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (audio_if_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (audio_if_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (audio_if_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (audio_if_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (audio_if_0_avalon_slave_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (audio_if_0_avalon_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (audio_if_0_avalon_slave_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (audio_if_0_avalon_slave_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (audio_if_0_avalon_slave_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (audio_if_0_avalon_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_007_source0_ready),                                                              //              cp.ready
		.cp_valid                (burst_adapter_007_source0_valid),                                                              //                .valid
		.cp_data                 (burst_adapter_007_source0_data),                                                               //                .data
		.cp_startofpacket        (burst_adapter_007_source0_startofpacket),                                                      //                .startofpacket
		.cp_endofpacket          (burst_adapter_007_source0_endofpacket),                                                        //                .endofpacket
		.cp_channel              (burst_adapter_007_source0_channel),                                                            //                .channel
		.rf_sink_ready           (audio_if_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (audio_if_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (audio_if_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (audio_if_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (audio_if_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (audio_if_0_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (audio_if_0_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (audio_if_0_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (audio_if_0_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (audio_if_0_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (audio_if_0_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (audio_if_0_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (audio_if_0_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (audio_if_0_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (audio_if_0_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (audio_if_0_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                                        //     (terminated)
		.m0_writeresponserequest (),                                                                                             //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                                          //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (114),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) audio_if_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (pll_audio_outclk0_clk),                                                                        //       clk.clk
		.reset             (rst_controller_003_reset_out_reset),                                                           // clk_reset.reset
		.in_data           (audio_if_0_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (audio_if_0_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (audio_if_0_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (audio_if_0_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (audio_if_0_avalon_slave_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (audio_if_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (audio_if_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (audio_if_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (audio_if_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (audio_if_0_avalon_slave_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                                        // (terminated)
		.csr_read          (1'b0),                                                                                         // (terminated)
		.csr_write         (1'b0),                                                                                         // (terminated)
		.csr_readdata      (),                                                                                             // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                         // (terminated)
		.almost_full_data  (),                                                                                             // (terminated)
		.almost_empty_data (),                                                                                             // (terminated)
		.in_empty          (1'b0),                                                                                         // (terminated)
		.out_empty         (),                                                                                             // (terminated)
		.in_error          (1'b0),                                                                                         // (terminated)
		.out_error         (),                                                                                             // (terminated)
		.in_channel        (1'b0),                                                                                         // (terminated)
		.out_channel       ()                                                                                              // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (34),
		.FIFO_DEPTH          (2),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (0),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) audio_if_0_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (pll_audio_outclk0_clk),                                                                  //       clk.clk
		.reset             (rst_controller_003_reset_out_reset),                                                     // clk_reset.reset
		.in_data           (audio_if_0_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (audio_if_0_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (audio_if_0_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (audio_if_0_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (audio_if_0_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (audio_if_0_avalon_slave_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                                  // (terminated)
		.csr_read          (1'b0),                                                                                   // (terminated)
		.csr_write         (1'b0),                                                                                   // (terminated)
		.csr_readdata      (),                                                                                       // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                                   // (terminated)
		.almost_full_data  (),                                                                                       // (terminated)
		.almost_empty_data (),                                                                                       // (terminated)
		.in_startofpacket  (1'b0),                                                                                   // (terminated)
		.in_endofpacket    (1'b0),                                                                                   // (terminated)
		.out_startofpacket (),                                                                                       // (terminated)
		.out_endofpacket   (),                                                                                       // (terminated)
		.in_empty          (1'b0),                                                                                   // (terminated)
		.out_empty         (),                                                                                       // (terminated)
		.in_error          (1'b0),                                                                                   // (terminated)
		.out_error         (),                                                                                       // (terminated)
		.in_channel        (1'b0),                                                                                   // (terminated)
		.out_channel       ()                                                                                        // (terminated)
	);

	altera_merlin_axi_master_ni #(
		.ID_WIDTH                  (12),
		.ADDR_WIDTH                (30),
		.RDATA_WIDTH               (128),
		.WDATA_WIDTH               (128),
		.ADDR_USER_WIDTH           (1),
		.DATA_USER_WIDTH           (1),
		.AXI_BURST_LENGTH_WIDTH    (4),
		.AXI_LOCK_WIDTH            (2),
		.AXI_VERSION               ("AXI3"),
		.WRITE_ISSUING_CAPABILITY  (8),
		.READ_ISSUING_CAPABILITY   (8),
		.PKT_BEGIN_BURST           (209),
		.PKT_CACHE_H               (231),
		.PKT_CACHE_L               (228),
		.PKT_ADDR_SIDEBAND_H       (207),
		.PKT_ADDR_SIDEBAND_L       (207),
		.PKT_PROTECTION_H          (227),
		.PKT_PROTECTION_L          (225),
		.PKT_BURST_SIZE_H          (204),
		.PKT_BURST_SIZE_L          (202),
		.PKT_BURST_TYPE_H          (206),
		.PKT_BURST_TYPE_L          (205),
		.PKT_RESPONSE_STATUS_L     (232),
		.PKT_RESPONSE_STATUS_H     (233),
		.PKT_BURSTWRAP_H           (201),
		.PKT_BURSTWRAP_L           (193),
		.PKT_BYTE_CNT_H            (192),
		.PKT_BYTE_CNT_L            (182),
		.PKT_ADDR_H                (175),
		.PKT_ADDR_L                (144),
		.PKT_TRANS_EXCLUSIVE       (181),
		.PKT_TRANS_LOCK            (180),
		.PKT_TRANS_COMPRESSED_READ (176),
		.PKT_TRANS_POSTED          (177),
		.PKT_TRANS_WRITE           (178),
		.PKT_TRANS_READ            (179),
		.PKT_DATA_H                (127),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (143),
		.PKT_BYTEEN_L              (128),
		.PKT_SRC_ID_H              (211),
		.PKT_SRC_ID_L              (211),
		.PKT_DEST_ID_H             (212),
		.PKT_DEST_ID_L             (212),
		.PKT_THREAD_ID_H           (224),
		.PKT_THREAD_ID_L           (213),
		.PKT_QOS_L                 (210),
		.PKT_QOS_H                 (210),
		.PKT_DATA_SIDEBAND_H       (208),
		.PKT_DATA_SIDEBAND_L       (208),
		.ST_DATA_W                 (234),
		.ST_CHANNEL_W              (3),
		.ID                        (1)
	) hps_0_h2f_axi_master_agent (
		.aclk                   (pll_sdram_outclk1_clk),                             //              clk.clk
		.aresetn                (~rst_controller_005_reset_out_reset),               //        clk_reset.reset_n
		.write_cp_valid         (hps_0_h2f_axi_master_agent_write_cp_valid),         //         write_cp.valid
		.write_cp_data          (hps_0_h2f_axi_master_agent_write_cp_data),          //                 .data
		.write_cp_startofpacket (hps_0_h2f_axi_master_agent_write_cp_startofpacket), //                 .startofpacket
		.write_cp_endofpacket   (hps_0_h2f_axi_master_agent_write_cp_endofpacket),   //                 .endofpacket
		.write_cp_ready         (hps_0_h2f_axi_master_agent_write_cp_ready),         //                 .ready
		.write_rp_valid         (rsp_xbar_demux_010_src0_valid),                     //         write_rp.valid
		.write_rp_data          (rsp_xbar_demux_010_src0_data),                      //                 .data
		.write_rp_channel       (rsp_xbar_demux_010_src0_channel),                   //                 .channel
		.write_rp_startofpacket (rsp_xbar_demux_010_src0_startofpacket),             //                 .startofpacket
		.write_rp_endofpacket   (rsp_xbar_demux_010_src0_endofpacket),               //                 .endofpacket
		.write_rp_ready         (rsp_xbar_demux_010_src0_ready),                     //                 .ready
		.read_cp_valid          (hps_0_h2f_axi_master_agent_read_cp_valid),          //          read_cp.valid
		.read_cp_data           (hps_0_h2f_axi_master_agent_read_cp_data),           //                 .data
		.read_cp_startofpacket  (hps_0_h2f_axi_master_agent_read_cp_startofpacket),  //                 .startofpacket
		.read_cp_endofpacket    (hps_0_h2f_axi_master_agent_read_cp_endofpacket),    //                 .endofpacket
		.read_cp_ready          (hps_0_h2f_axi_master_agent_read_cp_ready),          //                 .ready
		.read_rp_valid          (rsp_xbar_demux_010_src1_valid),                     //          read_rp.valid
		.read_rp_data           (rsp_xbar_demux_010_src1_data),                      //                 .data
		.read_rp_channel        (rsp_xbar_demux_010_src1_channel),                   //                 .channel
		.read_rp_startofpacket  (rsp_xbar_demux_010_src1_startofpacket),             //                 .startofpacket
		.read_rp_endofpacket    (rsp_xbar_demux_010_src1_endofpacket),               //                 .endofpacket
		.read_rp_ready          (rsp_xbar_demux_010_src1_ready),                     //                 .ready
		.awid                   (hps_0_h2f_axi_master_awid),                         // altera_axi_slave.awid
		.awaddr                 (hps_0_h2f_axi_master_awaddr),                       //                 .awaddr
		.awlen                  (hps_0_h2f_axi_master_awlen),                        //                 .awlen
		.awsize                 (hps_0_h2f_axi_master_awsize),                       //                 .awsize
		.awburst                (hps_0_h2f_axi_master_awburst),                      //                 .awburst
		.awlock                 (hps_0_h2f_axi_master_awlock),                       //                 .awlock
		.awcache                (hps_0_h2f_axi_master_awcache),                      //                 .awcache
		.awprot                 (hps_0_h2f_axi_master_awprot),                       //                 .awprot
		.awvalid                (hps_0_h2f_axi_master_awvalid),                      //                 .awvalid
		.awready                (hps_0_h2f_axi_master_awready),                      //                 .awready
		.wid                    (hps_0_h2f_axi_master_wid),                          //                 .wid
		.wdata                  (hps_0_h2f_axi_master_wdata),                        //                 .wdata
		.wstrb                  (hps_0_h2f_axi_master_wstrb),                        //                 .wstrb
		.wlast                  (hps_0_h2f_axi_master_wlast),                        //                 .wlast
		.wvalid                 (hps_0_h2f_axi_master_wvalid),                       //                 .wvalid
		.wready                 (hps_0_h2f_axi_master_wready),                       //                 .wready
		.bid                    (hps_0_h2f_axi_master_bid),                          //                 .bid
		.bresp                  (hps_0_h2f_axi_master_bresp),                        //                 .bresp
		.bvalid                 (hps_0_h2f_axi_master_bvalid),                       //                 .bvalid
		.bready                 (hps_0_h2f_axi_master_bready),                       //                 .bready
		.arid                   (hps_0_h2f_axi_master_arid),                         //                 .arid
		.araddr                 (hps_0_h2f_axi_master_araddr),                       //                 .araddr
		.arlen                  (hps_0_h2f_axi_master_arlen),                        //                 .arlen
		.arsize                 (hps_0_h2f_axi_master_arsize),                       //                 .arsize
		.arburst                (hps_0_h2f_axi_master_arburst),                      //                 .arburst
		.arlock                 (hps_0_h2f_axi_master_arlock),                       //                 .arlock
		.arcache                (hps_0_h2f_axi_master_arcache),                      //                 .arcache
		.arprot                 (hps_0_h2f_axi_master_arprot),                       //                 .arprot
		.arvalid                (hps_0_h2f_axi_master_arvalid),                      //                 .arvalid
		.arready                (hps_0_h2f_axi_master_arready),                      //                 .arready
		.rid                    (hps_0_h2f_axi_master_rid),                          //                 .rid
		.rdata                  (hps_0_h2f_axi_master_rdata),                        //                 .rdata
		.rresp                  (hps_0_h2f_axi_master_rresp),                        //                 .rresp
		.rlast                  (hps_0_h2f_axi_master_rlast),                        //                 .rlast
		.rvalid                 (hps_0_h2f_axi_master_rvalid),                       //                 .rvalid
		.rready                 (hps_0_h2f_axi_master_rready),                       //                 .rready
		.awuser                 (1'b0),                                              //      (terminated)
		.aruser                 (1'b0),                                              //      (terminated)
		.awqos                  (4'b0000),                                           //      (terminated)
		.arqos                  (4'b0000),                                           //      (terminated)
		.awregion               (4'b0000),                                           //      (terminated)
		.arregion               (4'b0000),                                           //      (terminated)
		.wuser                  (1'b0),                                              //      (terminated)
		.ruser                  (),                                                  //      (terminated)
		.buser                  ()                                                   //      (terminated)
	);

	altera_merlin_master_agent #(
		.PKT_PROTECTION_H          (119),
		.PKT_PROTECTION_L          (117),
		.PKT_BEGIN_BURST           (101),
		.PKT_BURSTWRAP_H           (93),
		.PKT_BURSTWRAP_L           (85),
		.PKT_BURST_SIZE_H          (96),
		.PKT_BURST_SIZE_L          (94),
		.PKT_BURST_TYPE_H          (98),
		.PKT_BURST_TYPE_L          (97),
		.PKT_BYTE_CNT_H            (84),
		.PKT_BYTE_CNT_L            (74),
		.PKT_ADDR_H                (67),
		.PKT_ADDR_L                (36),
		.PKT_TRANS_COMPRESSED_READ (68),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.PKT_TRANS_READ            (71),
		.PKT_TRANS_LOCK            (72),
		.PKT_TRANS_EXCLUSIVE       (73),
		.PKT_DATA_H                (31),
		.PKT_DATA_L                (0),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_SRC_ID_H              (103),
		.PKT_SRC_ID_L              (103),
		.PKT_DEST_ID_H             (104),
		.PKT_DEST_ID_L             (104),
		.PKT_THREAD_ID_H           (116),
		.PKT_THREAD_ID_L           (105),
		.PKT_CACHE_H               (123),
		.PKT_CACHE_L               (120),
		.PKT_DATA_SIDEBAND_H       (100),
		.PKT_DATA_SIDEBAND_L       (100),
		.PKT_QOS_H                 (102),
		.PKT_QOS_L                 (102),
		.PKT_ADDR_SIDEBAND_H       (99),
		.PKT_ADDR_SIDEBAND_L       (99),
		.PKT_RESPONSE_STATUS_H     (125),
		.PKT_RESPONSE_STATUS_L     (124),
		.ST_DATA_W                 (126),
		.ST_CHANNEL_W              (3),
		.AV_BURSTCOUNT_W           (9),
		.SUPPRESS_0_BYTEEN_RSP     (0),
		.ID                        (0),
		.BURSTWRAP_VALUE           (511),
		.CACHE_VALUE               (0),
		.SECURE_ACCESS_BIT         (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) alt_vip_vfr_0_avalon_master_translator_avalon_universal_master_0_agent (
		.clk                     (pll_sdram_outclk1_clk),                                                                   //       clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                                      // clk_reset.reset
		.av_address              (alt_vip_vfr_0_avalon_master_translator_avalon_universal_master_0_address),                //        av.address
		.av_write                (alt_vip_vfr_0_avalon_master_translator_avalon_universal_master_0_write),                  //          .write
		.av_read                 (alt_vip_vfr_0_avalon_master_translator_avalon_universal_master_0_read),                   //          .read
		.av_writedata            (alt_vip_vfr_0_avalon_master_translator_avalon_universal_master_0_writedata),              //          .writedata
		.av_readdata             (alt_vip_vfr_0_avalon_master_translator_avalon_universal_master_0_readdata),               //          .readdata
		.av_waitrequest          (alt_vip_vfr_0_avalon_master_translator_avalon_universal_master_0_waitrequest),            //          .waitrequest
		.av_readdatavalid        (alt_vip_vfr_0_avalon_master_translator_avalon_universal_master_0_readdatavalid),          //          .readdatavalid
		.av_byteenable           (alt_vip_vfr_0_avalon_master_translator_avalon_universal_master_0_byteenable),             //          .byteenable
		.av_burstcount           (alt_vip_vfr_0_avalon_master_translator_avalon_universal_master_0_burstcount),             //          .burstcount
		.av_debugaccess          (alt_vip_vfr_0_avalon_master_translator_avalon_universal_master_0_debugaccess),            //          .debugaccess
		.av_lock                 (alt_vip_vfr_0_avalon_master_translator_avalon_universal_master_0_lock),                   //          .lock
		.cp_valid                (alt_vip_vfr_0_avalon_master_translator_avalon_universal_master_0_agent_cp_valid),         //        cp.valid
		.cp_data                 (alt_vip_vfr_0_avalon_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.cp_startofpacket        (alt_vip_vfr_0_avalon_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.cp_endofpacket          (alt_vip_vfr_0_avalon_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.cp_ready                (alt_vip_vfr_0_avalon_master_translator_avalon_universal_master_0_agent_cp_ready),         //          .ready
		.rp_valid                (width_adapter_002_rsp_source_valid),                                                      //        rp.valid
		.rp_data                 (width_adapter_002_rsp_source_data),                                                       //          .data
		.rp_channel              (width_adapter_002_rsp_source_channel),                                                    //          .channel
		.rp_startofpacket        (width_adapter_002_rsp_source_startofpacket),                                              //          .startofpacket
		.rp_endofpacket          (width_adapter_002_rsp_source_endofpacket),                                                //          .endofpacket
		.rp_ready                (width_adapter_002_rsp_source_ready),                                                      //          .ready
		.av_response             (),                                                                                        // (terminated)
		.av_writeresponserequest (1'b0),                                                                                    // (terminated)
		.av_writeresponsevalid   ()                                                                                         // (terminated)
	);

	altera_merlin_slave_agent #(
		.PKT_DATA_H                (15),
		.PKT_DATA_L                (0),
		.PKT_BEGIN_BURST           (83),
		.PKT_SYMBOL_W              (8),
		.PKT_BYTEEN_H              (17),
		.PKT_BYTEEN_L              (16),
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (18),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_POSTED          (51),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.PKT_TRANS_LOCK            (54),
		.PKT_SRC_ID_H              (85),
		.PKT_SRC_ID_L              (85),
		.PKT_DEST_ID_H             (86),
		.PKT_DEST_ID_L             (86),
		.PKT_BURSTWRAP_H           (75),
		.PKT_BURSTWRAP_L           (67),
		.PKT_BYTE_CNT_H            (66),
		.PKT_BYTE_CNT_L            (56),
		.PKT_PROTECTION_H          (101),
		.PKT_PROTECTION_L          (99),
		.PKT_RESPONSE_STATUS_H     (107),
		.PKT_RESPONSE_STATUS_L     (106),
		.PKT_BURST_SIZE_H          (78),
		.PKT_BURST_SIZE_L          (76),
		.ST_CHANNEL_W              (3),
		.ST_DATA_W                 (108),
		.AVS_BURSTCOUNT_W          (2),
		.SUPPRESS_0_BYTEEN_CMD     (1),
		.PREVENT_FIFO_OVERFLOW     (1),
		.USE_READRESPONSE          (0),
		.USE_WRITERESPONSE         (0)
	) sdram_s1_translator_avalon_universal_slave_0_agent (
		.clk                     (pll_sdram_outclk1_clk),                                                         //             clk.clk
		.reset                   (rst_controller_001_reset_out_reset),                                            //       clk_reset.reset
		.m0_address              (sdram_s1_translator_avalon_universal_slave_0_agent_m0_address),                 //              m0.address
		.m0_burstcount           (sdram_s1_translator_avalon_universal_slave_0_agent_m0_burstcount),              //                .burstcount
		.m0_byteenable           (sdram_s1_translator_avalon_universal_slave_0_agent_m0_byteenable),              //                .byteenable
		.m0_debugaccess          (sdram_s1_translator_avalon_universal_slave_0_agent_m0_debugaccess),             //                .debugaccess
		.m0_lock                 (sdram_s1_translator_avalon_universal_slave_0_agent_m0_lock),                    //                .lock
		.m0_readdata             (sdram_s1_translator_avalon_universal_slave_0_agent_m0_readdata),                //                .readdata
		.m0_readdatavalid        (sdram_s1_translator_avalon_universal_slave_0_agent_m0_readdatavalid),           //                .readdatavalid
		.m0_read                 (sdram_s1_translator_avalon_universal_slave_0_agent_m0_read),                    //                .read
		.m0_waitrequest          (sdram_s1_translator_avalon_universal_slave_0_agent_m0_waitrequest),             //                .waitrequest
		.m0_writedata            (sdram_s1_translator_avalon_universal_slave_0_agent_m0_writedata),               //                .writedata
		.m0_write                (sdram_s1_translator_avalon_universal_slave_0_agent_m0_write),                   //                .write
		.rp_endofpacket          (sdram_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),             //              rp.endofpacket
		.rp_ready                (sdram_s1_translator_avalon_universal_slave_0_agent_rp_ready),                   //                .ready
		.rp_valid                (sdram_s1_translator_avalon_universal_slave_0_agent_rp_valid),                   //                .valid
		.rp_data                 (sdram_s1_translator_avalon_universal_slave_0_agent_rp_data),                    //                .data
		.rp_startofpacket        (sdram_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket),           //                .startofpacket
		.cp_ready                (burst_adapter_008_source0_ready),                                               //              cp.ready
		.cp_valid                (burst_adapter_008_source0_valid),                                               //                .valid
		.cp_data                 (burst_adapter_008_source0_data),                                                //                .data
		.cp_startofpacket        (burst_adapter_008_source0_startofpacket),                                       //                .startofpacket
		.cp_endofpacket          (burst_adapter_008_source0_endofpacket),                                         //                .endofpacket
		.cp_channel              (burst_adapter_008_source0_channel),                                             //                .channel
		.rf_sink_ready           (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //         rf_sink.ready
		.rf_sink_valid           (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //                .valid
		.rf_sink_startofpacket   (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //                .startofpacket
		.rf_sink_endofpacket     (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //                .endofpacket
		.rf_sink_data            (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //                .data
		.rf_source_ready         (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //       rf_source.ready
		.rf_source_valid         (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //                .valid
		.rf_source_startofpacket (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //                .startofpacket
		.rf_source_endofpacket   (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //                .endofpacket
		.rf_source_data          (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //                .data
		.rdata_fifo_sink_ready   (sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready),       // rdata_fifo_sink.ready
		.rdata_fifo_sink_valid   (sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid),       //                .valid
		.rdata_fifo_sink_data    (sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),        //                .data
		.rdata_fifo_src_ready    (sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready),       //  rdata_fifo_src.ready
		.rdata_fifo_src_valid    (sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid),       //                .valid
		.rdata_fifo_src_data     (sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),        //                .data
		.m0_response             (2'b00),                                                                         //     (terminated)
		.m0_writeresponserequest (),                                                                              //     (terminated)
		.m0_writeresponsevalid   (1'b0)                                                                           //     (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (109),
		.FIFO_DEPTH          (8),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (1),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (1),
		.USE_MEMORY_BLOCKS   (0),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo (
		.clk               (pll_sdram_outclk1_clk),                                                         //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                            // clk_reset.reset
		.in_data           (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_data),             //        in.data
		.in_valid          (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_valid),            //          .valid
		.in_ready          (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_ready),            //          .ready
		.in_startofpacket  (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_startofpacket),    //          .startofpacket
		.in_endofpacket    (sdram_s1_translator_avalon_universal_slave_0_agent_rf_source_endofpacket),      //          .endofpacket
		.out_data          (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_data),          //       out.data
		.out_valid         (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_valid),         //          .valid
		.out_ready         (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_ready),         //          .ready
		.out_startofpacket (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_startofpacket), //          .startofpacket
		.out_endofpacket   (sdram_s1_translator_avalon_universal_slave_0_agent_rsp_fifo_out_endofpacket),   //          .endofpacket
		.csr_address       (2'b00),                                                                         // (terminated)
		.csr_read          (1'b0),                                                                          // (terminated)
		.csr_write         (1'b0),                                                                          // (terminated)
		.csr_readdata      (),                                                                              // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                          // (terminated)
		.almost_full_data  (),                                                                              // (terminated)
		.almost_empty_data (),                                                                              // (terminated)
		.in_empty          (1'b0),                                                                          // (terminated)
		.out_empty         (),                                                                              // (terminated)
		.in_error          (1'b0),                                                                          // (terminated)
		.out_error         (),                                                                              // (terminated)
		.in_channel        (1'b0),                                                                          // (terminated)
		.out_channel       ()                                                                               // (terminated)
	);

	altera_avalon_sc_fifo #(
		.SYMBOLS_PER_BEAT    (1),
		.BITS_PER_SYMBOL     (18),
		.FIFO_DEPTH          (8),
		.CHANNEL_WIDTH       (0),
		.ERROR_WIDTH         (0),
		.USE_PACKETS         (0),
		.USE_FILL_LEVEL      (0),
		.EMPTY_LATENCY       (3),
		.USE_MEMORY_BLOCKS   (1),
		.USE_STORE_FORWARD   (0),
		.USE_ALMOST_FULL_IF  (0),
		.USE_ALMOST_EMPTY_IF (0)
	) sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo (
		.clk               (pll_sdram_outclk1_clk),                                                   //       clk.clk
		.reset             (rst_controller_001_reset_out_reset),                                      // clk_reset.reset
		.in_data           (sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_data),  //        in.data
		.in_valid          (sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_valid), //          .valid
		.in_ready          (sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_src_ready), //          .ready
		.out_data          (sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_data),  //       out.data
		.out_valid         (sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_valid), //          .valid
		.out_ready         (sdram_s1_translator_avalon_universal_slave_0_agent_rdata_fifo_out_ready), //          .ready
		.csr_address       (2'b00),                                                                   // (terminated)
		.csr_read          (1'b0),                                                                    // (terminated)
		.csr_write         (1'b0),                                                                    // (terminated)
		.csr_readdata      (),                                                                        // (terminated)
		.csr_writedata     (32'b00000000000000000000000000000000),                                    // (terminated)
		.almost_full_data  (),                                                                        // (terminated)
		.almost_empty_data (),                                                                        // (terminated)
		.in_startofpacket  (1'b0),                                                                    // (terminated)
		.in_endofpacket    (1'b0),                                                                    // (terminated)
		.out_startofpacket (),                                                                        // (terminated)
		.out_endofpacket   (),                                                                        // (terminated)
		.in_empty          (1'b0),                                                                    // (terminated)
		.out_empty         (),                                                                        // (terminated)
		.in_error          (1'b0),                                                                    // (terminated)
		.out_error         (),                                                                        // (terminated)
		.in_channel        (1'b0),                                                                    // (terminated)
		.out_channel       ()                                                                         // (terminated)
	);

	soc_system_addr_router addr_router (
		.sink_ready         (master_secure_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (master_secure_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (master_secure_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (master_secure_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (master_secure_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                          //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                   // clk_reset.reset
		.src_ready          (addr_router_src_ready),                                                            //       src.ready
		.src_valid          (addr_router_src_valid),                                                            //          .valid
		.src_data           (addr_router_src_data),                                                             //          .data
		.src_channel        (addr_router_src_channel),                                                          //          .channel
		.src_startofpacket  (addr_router_src_startofpacket),                                                    //          .startofpacket
		.src_endofpacket    (addr_router_src_endofpacket)                                                       //          .endofpacket
	);

	soc_system_id_router id_router (
		.sink_ready         (hps_0_f2h_axi_slave_agent_write_rp_ready),         //      sink.ready
		.sink_valid         (hps_0_f2h_axi_slave_agent_write_rp_valid),         //          .valid
		.sink_data          (hps_0_f2h_axi_slave_agent_write_rp_data),          //          .data
		.sink_startofpacket (hps_0_f2h_axi_slave_agent_write_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (hps_0_f2h_axi_slave_agent_write_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                          //       clk.clk
		.reset              (rst_controller_004_reset_out_reset),               // clk_reset.reset
		.src_ready          (id_router_src_ready),                              //       src.ready
		.src_valid          (id_router_src_valid),                              //          .valid
		.src_data           (id_router_src_data),                               //          .data
		.src_channel        (id_router_src_channel),                            //          .channel
		.src_startofpacket  (id_router_src_startofpacket),                      //          .startofpacket
		.src_endofpacket    (id_router_src_endofpacket)                         //          .endofpacket
	);

	soc_system_id_router id_router_001 (
		.sink_ready         (hps_0_f2h_axi_slave_agent_read_rp_ready),         //      sink.ready
		.sink_valid         (hps_0_f2h_axi_slave_agent_read_rp_valid),         //          .valid
		.sink_data          (hps_0_f2h_axi_slave_agent_read_rp_data),          //          .data
		.sink_startofpacket (hps_0_f2h_axi_slave_agent_read_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (hps_0_f2h_axi_slave_agent_read_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                         //       clk.clk
		.reset              (rst_controller_004_reset_out_reset),              // clk_reset.reset
		.src_ready          (id_router_001_src_ready),                         //       src.ready
		.src_valid          (id_router_001_src_valid),                         //          .valid
		.src_data           (id_router_001_src_data),                          //          .data
		.src_channel        (id_router_001_src_channel),                       //          .channel
		.src_startofpacket  (id_router_001_src_startofpacket),                 //          .startofpacket
		.src_endofpacket    (id_router_001_src_endofpacket)                    //          .endofpacket
	);

	soc_system_addr_router_001 addr_router_001 (
		.sink_ready         (hps_0_h2f_lw_axi_master_agent_write_cp_ready),         //      sink.ready
		.sink_valid         (hps_0_h2f_lw_axi_master_agent_write_cp_valid),         //          .valid
		.sink_data          (hps_0_h2f_lw_axi_master_agent_write_cp_data),          //          .data
		.sink_startofpacket (hps_0_h2f_lw_axi_master_agent_write_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (hps_0_h2f_lw_axi_master_agent_write_cp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                              //       clk.clk
		.reset              (rst_controller_004_reset_out_reset),                   // clk_reset.reset
		.src_ready          (addr_router_001_src_ready),                            //       src.ready
		.src_valid          (addr_router_001_src_valid),                            //          .valid
		.src_data           (addr_router_001_src_data),                             //          .data
		.src_channel        (addr_router_001_src_channel),                          //          .channel
		.src_startofpacket  (addr_router_001_src_startofpacket),                    //          .startofpacket
		.src_endofpacket    (addr_router_001_src_endofpacket)                       //          .endofpacket
	);

	soc_system_addr_router_001 addr_router_002 (
		.sink_ready         (hps_0_h2f_lw_axi_master_agent_read_cp_ready),         //      sink.ready
		.sink_valid         (hps_0_h2f_lw_axi_master_agent_read_cp_valid),         //          .valid
		.sink_data          (hps_0_h2f_lw_axi_master_agent_read_cp_data),          //          .data
		.sink_startofpacket (hps_0_h2f_lw_axi_master_agent_read_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (hps_0_h2f_lw_axi_master_agent_read_cp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                             //       clk.clk
		.reset              (rst_controller_004_reset_out_reset),                  // clk_reset.reset
		.src_ready          (addr_router_002_src_ready),                           //       src.ready
		.src_valid          (addr_router_002_src_valid),                           //          .valid
		.src_data           (addr_router_002_src_data),                            //          .data
		.src_channel        (addr_router_002_src_channel),                         //          .channel
		.src_startofpacket  (addr_router_002_src_startofpacket),                   //          .startofpacket
		.src_endofpacket    (addr_router_002_src_endofpacket)                      //          .endofpacket
	);

	soc_system_id_router_002 id_router_002 (
		.sink_ready         (led_pio_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (led_pio_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (led_pio_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (led_pio_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (led_pio_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                        // clk_reset.reset
		.src_ready          (id_router_002_src_ready),                                               //       src.ready
		.src_valid          (id_router_002_src_valid),                                               //          .valid
		.src_data           (id_router_002_src_data),                                                //          .data
		.src_channel        (id_router_002_src_channel),                                             //          .channel
		.src_startofpacket  (id_router_002_src_startofpacket),                                       //          .startofpacket
		.src_endofpacket    (id_router_002_src_endofpacket)                                          //          .endofpacket
	);

	soc_system_id_router_002 id_router_003 (
		.sink_ready         (dipsw_pio_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (dipsw_pio_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (dipsw_pio_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (dipsw_pio_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (dipsw_pio_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                 //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                          // clk_reset.reset
		.src_ready          (id_router_003_src_ready),                                                 //       src.ready
		.src_valid          (id_router_003_src_valid),                                                 //          .valid
		.src_data           (id_router_003_src_data),                                                  //          .data
		.src_channel        (id_router_003_src_channel),                                               //          .channel
		.src_startofpacket  (id_router_003_src_startofpacket),                                         //          .startofpacket
		.src_endofpacket    (id_router_003_src_endofpacket)                                            //          .endofpacket
	);

	soc_system_id_router_002 id_router_004 (
		.sink_ready         (button_pio_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (button_pio_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (button_pio_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (button_pio_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (button_pio_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                  //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                           // clk_reset.reset
		.src_ready          (id_router_004_src_ready),                                                  //       src.ready
		.src_valid          (id_router_004_src_valid),                                                  //          .valid
		.src_data           (id_router_004_src_data),                                                   //          .data
		.src_channel        (id_router_004_src_channel),                                                //          .channel
		.src_startofpacket  (id_router_004_src_startofpacket),                                          //          .startofpacket
		.src_endofpacket    (id_router_004_src_endofpacket)                                             //          .endofpacket
	);

	soc_system_id_router_002 id_router_005 (
		.sink_ready         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (jtag_uart_avalon_jtag_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                                //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                         // clk_reset.reset
		.src_ready          (id_router_005_src_ready),                                                                //       src.ready
		.src_valid          (id_router_005_src_valid),                                                                //          .valid
		.src_data           (id_router_005_src_data),                                                                 //          .data
		.src_channel        (id_router_005_src_channel),                                                              //          .channel
		.src_startofpacket  (id_router_005_src_startofpacket),                                                        //          .startofpacket
		.src_endofpacket    (id_router_005_src_endofpacket)                                                           //          .endofpacket
	);

	soc_system_id_router_002 id_router_006 (
		.sink_ready         (oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (oc_i2c_master_0_avalon_slave_0_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (clk_clk),                                                                                   //       clk.clk
		.reset              (rst_controller_reset_out_reset),                                                            // clk_reset.reset
		.src_ready          (id_router_006_src_ready),                                                                   //       src.ready
		.src_valid          (id_router_006_src_valid),                                                                   //          .valid
		.src_data           (id_router_006_src_data),                                                                    //          .data
		.src_channel        (id_router_006_src_channel),                                                                 //          .channel
		.src_startofpacket  (id_router_006_src_startofpacket),                                                           //          .startofpacket
		.src_endofpacket    (id_router_006_src_endofpacket)                                                              //          .endofpacket
	);

	soc_system_id_router_002 id_router_007 (
		.sink_ready         (alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (alt_vip_mix_0_control_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (pll_stream_outclk1_clk),                                                           //       clk.clk
		.reset              (rst_controller_002_reset_out_reset),                                               // clk_reset.reset
		.src_ready          (id_router_007_src_ready),                                                          //       src.ready
		.src_valid          (id_router_007_src_valid),                                                          //          .valid
		.src_data           (id_router_007_src_data),                                                           //          .data
		.src_channel        (id_router_007_src_channel),                                                        //          .channel
		.src_startofpacket  (id_router_007_src_startofpacket),                                                  //          .startofpacket
		.src_endofpacket    (id_router_007_src_endofpacket)                                                     //          .endofpacket
	);

	soc_system_id_router_002 id_router_008 (
		.sink_ready         (alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (alt_vip_vfr_0_avalon_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (pll_stream_outclk1_clk),                                                                //       clk.clk
		.reset              (rst_controller_002_reset_out_reset),                                                    // clk_reset.reset
		.src_ready          (id_router_008_src_ready),                                                               //       src.ready
		.src_valid          (id_router_008_src_valid),                                                               //          .valid
		.src_data           (id_router_008_src_data),                                                                //          .data
		.src_channel        (id_router_008_src_channel),                                                             //          .channel
		.src_startofpacket  (id_router_008_src_startofpacket),                                                       //          .startofpacket
		.src_endofpacket    (id_router_008_src_endofpacket)                                                          //          .endofpacket
	);

	soc_system_id_router_002 id_router_009 (
		.sink_ready         (audio_if_0_avalon_slave_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (audio_if_0_avalon_slave_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (audio_if_0_avalon_slave_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (audio_if_0_avalon_slave_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (audio_if_0_avalon_slave_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (pll_audio_outclk0_clk),                                                              //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),                                                 // clk_reset.reset
		.src_ready          (id_router_009_src_ready),                                                            //       src.ready
		.src_valid          (id_router_009_src_valid),                                                            //          .valid
		.src_data           (id_router_009_src_data),                                                             //          .data
		.src_channel        (id_router_009_src_channel),                                                          //          .channel
		.src_startofpacket  (id_router_009_src_startofpacket),                                                    //          .startofpacket
		.src_endofpacket    (id_router_009_src_endofpacket)                                                       //          .endofpacket
	);

	soc_system_addr_router_003 addr_router_003 (
		.sink_ready         (hps_0_h2f_axi_master_agent_write_cp_ready),         //      sink.ready
		.sink_valid         (hps_0_h2f_axi_master_agent_write_cp_valid),         //          .valid
		.sink_data          (hps_0_h2f_axi_master_agent_write_cp_data),          //          .data
		.sink_startofpacket (hps_0_h2f_axi_master_agent_write_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (hps_0_h2f_axi_master_agent_write_cp_endofpacket),   //          .endofpacket
		.clk                (pll_sdram_outclk1_clk),                             //       clk.clk
		.reset              (rst_controller_005_reset_out_reset),                // clk_reset.reset
		.src_ready          (addr_router_003_src_ready),                         //       src.ready
		.src_valid          (addr_router_003_src_valid),                         //          .valid
		.src_data           (addr_router_003_src_data),                          //          .data
		.src_channel        (addr_router_003_src_channel),                       //          .channel
		.src_startofpacket  (addr_router_003_src_startofpacket),                 //          .startofpacket
		.src_endofpacket    (addr_router_003_src_endofpacket)                    //          .endofpacket
	);

	soc_system_addr_router_003 addr_router_004 (
		.sink_ready         (hps_0_h2f_axi_master_agent_read_cp_ready),         //      sink.ready
		.sink_valid         (hps_0_h2f_axi_master_agent_read_cp_valid),         //          .valid
		.sink_data          (hps_0_h2f_axi_master_agent_read_cp_data),          //          .data
		.sink_startofpacket (hps_0_h2f_axi_master_agent_read_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (hps_0_h2f_axi_master_agent_read_cp_endofpacket),   //          .endofpacket
		.clk                (pll_sdram_outclk1_clk),                            //       clk.clk
		.reset              (rst_controller_005_reset_out_reset),               // clk_reset.reset
		.src_ready          (addr_router_004_src_ready),                        //       src.ready
		.src_valid          (addr_router_004_src_valid),                        //          .valid
		.src_data           (addr_router_004_src_data),                         //          .data
		.src_channel        (addr_router_004_src_channel),                      //          .channel
		.src_startofpacket  (addr_router_004_src_startofpacket),                //          .startofpacket
		.src_endofpacket    (addr_router_004_src_endofpacket)                   //          .endofpacket
	);

	soc_system_addr_router_005 addr_router_005 (
		.sink_ready         (alt_vip_vfr_0_avalon_master_translator_avalon_universal_master_0_agent_cp_ready),         //      sink.ready
		.sink_valid         (alt_vip_vfr_0_avalon_master_translator_avalon_universal_master_0_agent_cp_valid),         //          .valid
		.sink_data          (alt_vip_vfr_0_avalon_master_translator_avalon_universal_master_0_agent_cp_data),          //          .data
		.sink_startofpacket (alt_vip_vfr_0_avalon_master_translator_avalon_universal_master_0_agent_cp_startofpacket), //          .startofpacket
		.sink_endofpacket   (alt_vip_vfr_0_avalon_master_translator_avalon_universal_master_0_agent_cp_endofpacket),   //          .endofpacket
		.clk                (pll_sdram_outclk1_clk),                                                                   //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                                      // clk_reset.reset
		.src_ready          (addr_router_005_src_ready),                                                               //       src.ready
		.src_valid          (addr_router_005_src_valid),                                                               //          .valid
		.src_data           (addr_router_005_src_data),                                                                //          .data
		.src_channel        (addr_router_005_src_channel),                                                             //          .channel
		.src_startofpacket  (addr_router_005_src_startofpacket),                                                       //          .startofpacket
		.src_endofpacket    (addr_router_005_src_endofpacket)                                                          //          .endofpacket
	);

	soc_system_id_router_010 id_router_010 (
		.sink_ready         (sdram_s1_translator_avalon_universal_slave_0_agent_rp_ready),         //      sink.ready
		.sink_valid         (sdram_s1_translator_avalon_universal_slave_0_agent_rp_valid),         //          .valid
		.sink_data          (sdram_s1_translator_avalon_universal_slave_0_agent_rp_data),          //          .data
		.sink_startofpacket (sdram_s1_translator_avalon_universal_slave_0_agent_rp_startofpacket), //          .startofpacket
		.sink_endofpacket   (sdram_s1_translator_avalon_universal_slave_0_agent_rp_endofpacket),   //          .endofpacket
		.clk                (pll_sdram_outclk1_clk),                                               //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),                                  // clk_reset.reset
		.src_ready          (id_router_010_src_ready),                                             //       src.ready
		.src_valid          (id_router_010_src_valid),                                             //          .valid
		.src_data           (id_router_010_src_data),                                              //          .data
		.src_channel        (id_router_010_src_channel),                                           //          .channel
		.src_startofpacket  (id_router_010_src_startofpacket),                                     //          .startofpacket
		.src_endofpacket    (id_router_010_src_endofpacket)                                        //          .endofpacket
	);

	altera_merlin_traffic_limiter #(
		.PKT_DEST_ID_H             (104),
		.PKT_DEST_ID_L             (104),
		.PKT_TRANS_POSTED          (69),
		.PKT_TRANS_WRITE           (70),
		.MAX_OUTSTANDING_RESPONSES (16),
		.PIPELINED                 (0),
		.ST_DATA_W                 (115),
		.ST_CHANNEL_W              (2),
		.VALID_WIDTH               (2),
		.ENFORCE_ORDER             (1),
		.PREVENT_HAZARDS           (1),
		.PKT_BYTE_CNT_H            (81),
		.PKT_BYTE_CNT_L            (74),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32)
	) limiter (
		.clk                    (clk_clk),                        //       clk.clk
		.reset                  (rst_controller_reset_out_reset), // clk_reset.reset
		.cmd_sink_ready         (addr_router_src_ready),          //  cmd_sink.ready
		.cmd_sink_valid         (addr_router_src_valid),          //          .valid
		.cmd_sink_data          (addr_router_src_data),           //          .data
		.cmd_sink_channel       (addr_router_src_channel),        //          .channel
		.cmd_sink_startofpacket (addr_router_src_startofpacket),  //          .startofpacket
		.cmd_sink_endofpacket   (addr_router_src_endofpacket),    //          .endofpacket
		.cmd_src_ready          (limiter_cmd_src_ready),          //   cmd_src.ready
		.cmd_src_data           (limiter_cmd_src_data),           //          .data
		.cmd_src_channel        (limiter_cmd_src_channel),        //          .channel
		.cmd_src_startofpacket  (limiter_cmd_src_startofpacket),  //          .startofpacket
		.cmd_src_endofpacket    (limiter_cmd_src_endofpacket),    //          .endofpacket
		.rsp_sink_ready         (rsp_xbar_mux_src_ready),         //  rsp_sink.ready
		.rsp_sink_valid         (rsp_xbar_mux_src_valid),         //          .valid
		.rsp_sink_channel       (rsp_xbar_mux_src_channel),       //          .channel
		.rsp_sink_data          (rsp_xbar_mux_src_data),          //          .data
		.rsp_sink_startofpacket (rsp_xbar_mux_src_startofpacket), //          .startofpacket
		.rsp_sink_endofpacket   (rsp_xbar_mux_src_endofpacket),   //          .endofpacket
		.rsp_src_ready          (limiter_rsp_src_ready),          //   rsp_src.ready
		.rsp_src_valid          (limiter_rsp_src_valid),          //          .valid
		.rsp_src_data           (limiter_rsp_src_data),           //          .data
		.rsp_src_channel        (limiter_rsp_src_channel),        //          .channel
		.rsp_src_startofpacket  (limiter_rsp_src_startofpacket),  //          .startofpacket
		.rsp_src_endofpacket    (limiter_rsp_src_endofpacket),    //          .endofpacket
		.cmd_src_valid          (limiter_cmd_valid_data)          // cmd_valid.data
	);

	altera_merlin_traffic_limiter #(
		.PKT_DEST_ID_H             (91),
		.PKT_DEST_ID_L             (89),
		.PKT_TRANS_POSTED          (58),
		.PKT_TRANS_WRITE           (59),
		.MAX_OUTSTANDING_RESPONSES (7),
		.PIPELINED                 (0),
		.ST_DATA_W                 (113),
		.ST_CHANNEL_W              (8),
		.VALID_WIDTH               (8),
		.ENFORCE_ORDER             (1),
		.PREVENT_HAZARDS           (0),
		.PKT_BYTE_CNT_H            (69),
		.PKT_BYTE_CNT_L            (63),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32)
	) limiter_001 (
		.clk                    (clk_clk),                            //       clk.clk
		.reset                  (rst_controller_004_reset_out_reset), // clk_reset.reset
		.cmd_sink_ready         (addr_router_001_src_ready),          //  cmd_sink.ready
		.cmd_sink_valid         (addr_router_001_src_valid),          //          .valid
		.cmd_sink_data          (addr_router_001_src_data),           //          .data
		.cmd_sink_channel       (addr_router_001_src_channel),        //          .channel
		.cmd_sink_startofpacket (addr_router_001_src_startofpacket),  //          .startofpacket
		.cmd_sink_endofpacket   (addr_router_001_src_endofpacket),    //          .endofpacket
		.cmd_src_ready          (limiter_001_cmd_src_ready),          //   cmd_src.ready
		.cmd_src_data           (limiter_001_cmd_src_data),           //          .data
		.cmd_src_channel        (limiter_001_cmd_src_channel),        //          .channel
		.cmd_src_startofpacket  (limiter_001_cmd_src_startofpacket),  //          .startofpacket
		.cmd_src_endofpacket    (limiter_001_cmd_src_endofpacket),    //          .endofpacket
		.rsp_sink_ready         (rsp_xbar_mux_001_src_ready),         //  rsp_sink.ready
		.rsp_sink_valid         (rsp_xbar_mux_001_src_valid),         //          .valid
		.rsp_sink_channel       (rsp_xbar_mux_001_src_channel),       //          .channel
		.rsp_sink_data          (rsp_xbar_mux_001_src_data),          //          .data
		.rsp_sink_startofpacket (rsp_xbar_mux_001_src_startofpacket), //          .startofpacket
		.rsp_sink_endofpacket   (rsp_xbar_mux_001_src_endofpacket),   //          .endofpacket
		.rsp_src_ready          (limiter_001_rsp_src_ready),          //   rsp_src.ready
		.rsp_src_valid          (limiter_001_rsp_src_valid),          //          .valid
		.rsp_src_data           (limiter_001_rsp_src_data),           //          .data
		.rsp_src_channel        (limiter_001_rsp_src_channel),        //          .channel
		.rsp_src_startofpacket  (limiter_001_rsp_src_startofpacket),  //          .startofpacket
		.rsp_src_endofpacket    (limiter_001_rsp_src_endofpacket),    //          .endofpacket
		.cmd_src_valid          (limiter_001_cmd_valid_data)          // cmd_valid.data
	);

	altera_merlin_traffic_limiter #(
		.PKT_DEST_ID_H             (91),
		.PKT_DEST_ID_L             (89),
		.PKT_TRANS_POSTED          (58),
		.PKT_TRANS_WRITE           (59),
		.MAX_OUTSTANDING_RESPONSES (7),
		.PIPELINED                 (0),
		.ST_DATA_W                 (113),
		.ST_CHANNEL_W              (8),
		.VALID_WIDTH               (8),
		.ENFORCE_ORDER             (1),
		.PREVENT_HAZARDS           (0),
		.PKT_BYTE_CNT_H            (69),
		.PKT_BYTE_CNT_L            (63),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32)
	) limiter_002 (
		.clk                    (clk_clk),                            //       clk.clk
		.reset                  (rst_controller_004_reset_out_reset), // clk_reset.reset
		.cmd_sink_ready         (addr_router_002_src_ready),          //  cmd_sink.ready
		.cmd_sink_valid         (addr_router_002_src_valid),          //          .valid
		.cmd_sink_data          (addr_router_002_src_data),           //          .data
		.cmd_sink_channel       (addr_router_002_src_channel),        //          .channel
		.cmd_sink_startofpacket (addr_router_002_src_startofpacket),  //          .startofpacket
		.cmd_sink_endofpacket   (addr_router_002_src_endofpacket),    //          .endofpacket
		.cmd_src_ready          (limiter_002_cmd_src_ready),          //   cmd_src.ready
		.cmd_src_data           (limiter_002_cmd_src_data),           //          .data
		.cmd_src_channel        (limiter_002_cmd_src_channel),        //          .channel
		.cmd_src_startofpacket  (limiter_002_cmd_src_startofpacket),  //          .startofpacket
		.cmd_src_endofpacket    (limiter_002_cmd_src_endofpacket),    //          .endofpacket
		.rsp_sink_ready         (rsp_xbar_mux_002_src_ready),         //  rsp_sink.ready
		.rsp_sink_valid         (rsp_xbar_mux_002_src_valid),         //          .valid
		.rsp_sink_channel       (rsp_xbar_mux_002_src_channel),       //          .channel
		.rsp_sink_data          (rsp_xbar_mux_002_src_data),          //          .data
		.rsp_sink_startofpacket (rsp_xbar_mux_002_src_startofpacket), //          .startofpacket
		.rsp_sink_endofpacket   (rsp_xbar_mux_002_src_endofpacket),   //          .endofpacket
		.rsp_src_ready          (limiter_002_rsp_src_ready),          //   rsp_src.ready
		.rsp_src_valid          (limiter_002_rsp_src_valid),          //          .valid
		.rsp_src_data           (limiter_002_rsp_src_data),           //          .data
		.rsp_src_channel        (limiter_002_rsp_src_channel),        //          .channel
		.rsp_src_startofpacket  (limiter_002_rsp_src_startofpacket),  //          .startofpacket
		.rsp_src_endofpacket    (limiter_002_rsp_src_endofpacket),    //          .endofpacket
		.cmd_src_valid          (limiter_002_cmd_valid_data)          // cmd_valid.data
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (56),
		.PKT_ADDR_L                (36),
		.PKT_BEGIN_BURST           (84),
		.PKT_BYTE_CNT_H            (69),
		.PKT_BYTE_CNT_L            (63),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_BURST_SIZE_H          (79),
		.PKT_BURST_SIZE_L          (77),
		.PKT_BURST_TYPE_H          (81),
		.PKT_BURST_TYPE_L          (80),
		.PKT_BURSTWRAP_H           (76),
		.PKT_BURSTWRAP_L           (70),
		.PKT_TRANS_COMPRESSED_READ (57),
		.PKT_TRANS_WRITE           (59),
		.PKT_TRANS_READ            (60),
		.OUT_NARROW_SIZE           (0),
		.IN_NARROW_SIZE            (1),
		.OUT_FIXED                 (0),
		.OUT_COMPLETE_WRAP         (0),
		.ST_DATA_W                 (113),
		.ST_CHANNEL_W              (8),
		.OUT_BYTE_CNT_H            (65),
		.OUT_BURSTWRAP_H           (76),
		.COMPRESSED_READ_SUPPORT   (1),
		.BYTEENABLE_SYNTHESIS      (1),
		.PIPE_INPUTS               (0),
		.NO_WRAP_SUPPORT           (0),
		.BURSTWRAP_CONST_MASK      (0),
		.BURSTWRAP_CONST_VALUE     (0)
	) burst_adapter (
		.clk                   (clk_clk),                             //       cr0.clk
		.reset                 (rst_controller_reset_out_reset),      // cr0_reset.reset
		.sink0_valid           (cmd_xbar_mux_002_src_valid),          //     sink0.valid
		.sink0_data            (cmd_xbar_mux_002_src_data),           //          .data
		.sink0_channel         (cmd_xbar_mux_002_src_channel),        //          .channel
		.sink0_startofpacket   (cmd_xbar_mux_002_src_startofpacket),  //          .startofpacket
		.sink0_endofpacket     (cmd_xbar_mux_002_src_endofpacket),    //          .endofpacket
		.sink0_ready           (cmd_xbar_mux_002_src_ready),          //          .ready
		.source0_valid         (burst_adapter_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_source0_data),          //          .data
		.source0_channel       (burst_adapter_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_source0_ready)          //          .ready
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (56),
		.PKT_ADDR_L                (36),
		.PKT_BEGIN_BURST           (84),
		.PKT_BYTE_CNT_H            (69),
		.PKT_BYTE_CNT_L            (63),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_BURST_SIZE_H          (79),
		.PKT_BURST_SIZE_L          (77),
		.PKT_BURST_TYPE_H          (81),
		.PKT_BURST_TYPE_L          (80),
		.PKT_BURSTWRAP_H           (76),
		.PKT_BURSTWRAP_L           (70),
		.PKT_TRANS_COMPRESSED_READ (57),
		.PKT_TRANS_WRITE           (59),
		.PKT_TRANS_READ            (60),
		.OUT_NARROW_SIZE           (0),
		.IN_NARROW_SIZE            (1),
		.OUT_FIXED                 (0),
		.OUT_COMPLETE_WRAP         (0),
		.ST_DATA_W                 (113),
		.ST_CHANNEL_W              (8),
		.OUT_BYTE_CNT_H            (65),
		.OUT_BURSTWRAP_H           (76),
		.COMPRESSED_READ_SUPPORT   (1),
		.BYTEENABLE_SYNTHESIS      (1),
		.PIPE_INPUTS               (0),
		.NO_WRAP_SUPPORT           (0),
		.BURSTWRAP_CONST_MASK      (0),
		.BURSTWRAP_CONST_VALUE     (0)
	) burst_adapter_001 (
		.clk                   (clk_clk),                                 //       cr0.clk
		.reset                 (rst_controller_reset_out_reset),          // cr0_reset.reset
		.sink0_valid           (cmd_xbar_mux_003_src_valid),              //     sink0.valid
		.sink0_data            (cmd_xbar_mux_003_src_data),               //          .data
		.sink0_channel         (cmd_xbar_mux_003_src_channel),            //          .channel
		.sink0_startofpacket   (cmd_xbar_mux_003_src_startofpacket),      //          .startofpacket
		.sink0_endofpacket     (cmd_xbar_mux_003_src_endofpacket),        //          .endofpacket
		.sink0_ready           (cmd_xbar_mux_003_src_ready),              //          .ready
		.source0_valid         (burst_adapter_001_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_001_source0_data),          //          .data
		.source0_channel       (burst_adapter_001_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_001_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_001_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_001_source0_ready)          //          .ready
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (56),
		.PKT_ADDR_L                (36),
		.PKT_BEGIN_BURST           (84),
		.PKT_BYTE_CNT_H            (69),
		.PKT_BYTE_CNT_L            (63),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_BURST_SIZE_H          (79),
		.PKT_BURST_SIZE_L          (77),
		.PKT_BURST_TYPE_H          (81),
		.PKT_BURST_TYPE_L          (80),
		.PKT_BURSTWRAP_H           (76),
		.PKT_BURSTWRAP_L           (70),
		.PKT_TRANS_COMPRESSED_READ (57),
		.PKT_TRANS_WRITE           (59),
		.PKT_TRANS_READ            (60),
		.OUT_NARROW_SIZE           (0),
		.IN_NARROW_SIZE            (1),
		.OUT_FIXED                 (0),
		.OUT_COMPLETE_WRAP         (0),
		.ST_DATA_W                 (113),
		.ST_CHANNEL_W              (8),
		.OUT_BYTE_CNT_H            (65),
		.OUT_BURSTWRAP_H           (76),
		.COMPRESSED_READ_SUPPORT   (1),
		.BYTEENABLE_SYNTHESIS      (1),
		.PIPE_INPUTS               (0),
		.NO_WRAP_SUPPORT           (0),
		.BURSTWRAP_CONST_MASK      (0),
		.BURSTWRAP_CONST_VALUE     (0)
	) burst_adapter_002 (
		.clk                   (clk_clk),                                 //       cr0.clk
		.reset                 (rst_controller_reset_out_reset),          // cr0_reset.reset
		.sink0_valid           (cmd_xbar_mux_004_src_valid),              //     sink0.valid
		.sink0_data            (cmd_xbar_mux_004_src_data),               //          .data
		.sink0_channel         (cmd_xbar_mux_004_src_channel),            //          .channel
		.sink0_startofpacket   (cmd_xbar_mux_004_src_startofpacket),      //          .startofpacket
		.sink0_endofpacket     (cmd_xbar_mux_004_src_endofpacket),        //          .endofpacket
		.sink0_ready           (cmd_xbar_mux_004_src_ready),              //          .ready
		.source0_valid         (burst_adapter_002_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_002_source0_data),          //          .data
		.source0_channel       (burst_adapter_002_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_002_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_002_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_002_source0_ready)          //          .ready
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (56),
		.PKT_ADDR_L                (36),
		.PKT_BEGIN_BURST           (84),
		.PKT_BYTE_CNT_H            (69),
		.PKT_BYTE_CNT_L            (63),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_BURST_SIZE_H          (79),
		.PKT_BURST_SIZE_L          (77),
		.PKT_BURST_TYPE_H          (81),
		.PKT_BURST_TYPE_L          (80),
		.PKT_BURSTWRAP_H           (76),
		.PKT_BURSTWRAP_L           (70),
		.PKT_TRANS_COMPRESSED_READ (57),
		.PKT_TRANS_WRITE           (59),
		.PKT_TRANS_READ            (60),
		.OUT_NARROW_SIZE           (0),
		.IN_NARROW_SIZE            (1),
		.OUT_FIXED                 (0),
		.OUT_COMPLETE_WRAP         (0),
		.ST_DATA_W                 (113),
		.ST_CHANNEL_W              (8),
		.OUT_BYTE_CNT_H            (65),
		.OUT_BURSTWRAP_H           (76),
		.COMPRESSED_READ_SUPPORT   (1),
		.BYTEENABLE_SYNTHESIS      (1),
		.PIPE_INPUTS               (0),
		.NO_WRAP_SUPPORT           (0),
		.BURSTWRAP_CONST_MASK      (0),
		.BURSTWRAP_CONST_VALUE     (0)
	) burst_adapter_003 (
		.clk                   (clk_clk),                                 //       cr0.clk
		.reset                 (rst_controller_reset_out_reset),          // cr0_reset.reset
		.sink0_valid           (cmd_xbar_mux_005_src_valid),              //     sink0.valid
		.sink0_data            (cmd_xbar_mux_005_src_data),               //          .data
		.sink0_channel         (cmd_xbar_mux_005_src_channel),            //          .channel
		.sink0_startofpacket   (cmd_xbar_mux_005_src_startofpacket),      //          .startofpacket
		.sink0_endofpacket     (cmd_xbar_mux_005_src_endofpacket),        //          .endofpacket
		.sink0_ready           (cmd_xbar_mux_005_src_ready),              //          .ready
		.source0_valid         (burst_adapter_003_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_003_source0_data),          //          .data
		.source0_channel       (burst_adapter_003_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_003_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_003_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_003_source0_ready)          //          .ready
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (56),
		.PKT_ADDR_L                (36),
		.PKT_BEGIN_BURST           (84),
		.PKT_BYTE_CNT_H            (69),
		.PKT_BYTE_CNT_L            (63),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_BURST_SIZE_H          (79),
		.PKT_BURST_SIZE_L          (77),
		.PKT_BURST_TYPE_H          (81),
		.PKT_BURST_TYPE_L          (80),
		.PKT_BURSTWRAP_H           (76),
		.PKT_BURSTWRAP_L           (70),
		.PKT_TRANS_COMPRESSED_READ (57),
		.PKT_TRANS_WRITE           (59),
		.PKT_TRANS_READ            (60),
		.OUT_NARROW_SIZE           (0),
		.IN_NARROW_SIZE            (1),
		.OUT_FIXED                 (0),
		.OUT_COMPLETE_WRAP         (0),
		.ST_DATA_W                 (113),
		.ST_CHANNEL_W              (8),
		.OUT_BYTE_CNT_H            (65),
		.OUT_BURSTWRAP_H           (76),
		.COMPRESSED_READ_SUPPORT   (1),
		.BYTEENABLE_SYNTHESIS      (1),
		.PIPE_INPUTS               (0),
		.NO_WRAP_SUPPORT           (0),
		.BURSTWRAP_CONST_MASK      (0),
		.BURSTWRAP_CONST_VALUE     (0)
	) burst_adapter_004 (
		.clk                   (clk_clk),                                 //       cr0.clk
		.reset                 (rst_controller_reset_out_reset),          // cr0_reset.reset
		.sink0_valid           (cmd_xbar_mux_006_src_valid),              //     sink0.valid
		.sink0_data            (cmd_xbar_mux_006_src_data),               //          .data
		.sink0_channel         (cmd_xbar_mux_006_src_channel),            //          .channel
		.sink0_startofpacket   (cmd_xbar_mux_006_src_startofpacket),      //          .startofpacket
		.sink0_endofpacket     (cmd_xbar_mux_006_src_endofpacket),        //          .endofpacket
		.sink0_ready           (cmd_xbar_mux_006_src_ready),              //          .ready
		.source0_valid         (burst_adapter_004_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_004_source0_data),          //          .data
		.source0_channel       (burst_adapter_004_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_004_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_004_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_004_source0_ready)          //          .ready
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (56),
		.PKT_ADDR_L                (36),
		.PKT_BEGIN_BURST           (84),
		.PKT_BYTE_CNT_H            (69),
		.PKT_BYTE_CNT_L            (63),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_BURST_SIZE_H          (79),
		.PKT_BURST_SIZE_L          (77),
		.PKT_BURST_TYPE_H          (81),
		.PKT_BURST_TYPE_L          (80),
		.PKT_BURSTWRAP_H           (76),
		.PKT_BURSTWRAP_L           (70),
		.PKT_TRANS_COMPRESSED_READ (57),
		.PKT_TRANS_WRITE           (59),
		.PKT_TRANS_READ            (60),
		.OUT_NARROW_SIZE           (0),
		.IN_NARROW_SIZE            (1),
		.OUT_FIXED                 (0),
		.OUT_COMPLETE_WRAP         (0),
		.ST_DATA_W                 (113),
		.ST_CHANNEL_W              (8),
		.OUT_BYTE_CNT_H            (65),
		.OUT_BURSTWRAP_H           (76),
		.COMPRESSED_READ_SUPPORT   (1),
		.BYTEENABLE_SYNTHESIS      (1),
		.PIPE_INPUTS               (0),
		.NO_WRAP_SUPPORT           (0),
		.BURSTWRAP_CONST_MASK      (0),
		.BURSTWRAP_CONST_VALUE     (0)
	) burst_adapter_005 (
		.clk                   (pll_stream_outclk1_clk),                  //       cr0.clk
		.reset                 (rst_controller_002_reset_out_reset),      // cr0_reset.reset
		.sink0_valid           (cmd_xbar_mux_007_src_valid),              //     sink0.valid
		.sink0_data            (cmd_xbar_mux_007_src_data),               //          .data
		.sink0_channel         (cmd_xbar_mux_007_src_channel),            //          .channel
		.sink0_startofpacket   (cmd_xbar_mux_007_src_startofpacket),      //          .startofpacket
		.sink0_endofpacket     (cmd_xbar_mux_007_src_endofpacket),        //          .endofpacket
		.sink0_ready           (cmd_xbar_mux_007_src_ready),              //          .ready
		.source0_valid         (burst_adapter_005_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_005_source0_data),          //          .data
		.source0_channel       (burst_adapter_005_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_005_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_005_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_005_source0_ready)          //          .ready
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (56),
		.PKT_ADDR_L                (36),
		.PKT_BEGIN_BURST           (84),
		.PKT_BYTE_CNT_H            (69),
		.PKT_BYTE_CNT_L            (63),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_BURST_SIZE_H          (79),
		.PKT_BURST_SIZE_L          (77),
		.PKT_BURST_TYPE_H          (81),
		.PKT_BURST_TYPE_L          (80),
		.PKT_BURSTWRAP_H           (76),
		.PKT_BURSTWRAP_L           (70),
		.PKT_TRANS_COMPRESSED_READ (57),
		.PKT_TRANS_WRITE           (59),
		.PKT_TRANS_READ            (60),
		.OUT_NARROW_SIZE           (0),
		.IN_NARROW_SIZE            (1),
		.OUT_FIXED                 (0),
		.OUT_COMPLETE_WRAP         (0),
		.ST_DATA_W                 (113),
		.ST_CHANNEL_W              (8),
		.OUT_BYTE_CNT_H            (65),
		.OUT_BURSTWRAP_H           (76),
		.COMPRESSED_READ_SUPPORT   (1),
		.BYTEENABLE_SYNTHESIS      (1),
		.PIPE_INPUTS               (0),
		.NO_WRAP_SUPPORT           (0),
		.BURSTWRAP_CONST_MASK      (0),
		.BURSTWRAP_CONST_VALUE     (0)
	) burst_adapter_006 (
		.clk                   (pll_stream_outclk1_clk),                  //       cr0.clk
		.reset                 (rst_controller_002_reset_out_reset),      // cr0_reset.reset
		.sink0_valid           (cmd_xbar_mux_008_src_valid),              //     sink0.valid
		.sink0_data            (cmd_xbar_mux_008_src_data),               //          .data
		.sink0_channel         (cmd_xbar_mux_008_src_channel),            //          .channel
		.sink0_startofpacket   (cmd_xbar_mux_008_src_startofpacket),      //          .startofpacket
		.sink0_endofpacket     (cmd_xbar_mux_008_src_endofpacket),        //          .endofpacket
		.sink0_ready           (cmd_xbar_mux_008_src_ready),              //          .ready
		.source0_valid         (burst_adapter_006_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_006_source0_data),          //          .data
		.source0_channel       (burst_adapter_006_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_006_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_006_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_006_source0_ready)          //          .ready
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (56),
		.PKT_ADDR_L                (36),
		.PKT_BEGIN_BURST           (84),
		.PKT_BYTE_CNT_H            (69),
		.PKT_BYTE_CNT_L            (63),
		.PKT_BYTEEN_H              (35),
		.PKT_BYTEEN_L              (32),
		.PKT_BURST_SIZE_H          (79),
		.PKT_BURST_SIZE_L          (77),
		.PKT_BURST_TYPE_H          (81),
		.PKT_BURST_TYPE_L          (80),
		.PKT_BURSTWRAP_H           (76),
		.PKT_BURSTWRAP_L           (70),
		.PKT_TRANS_COMPRESSED_READ (57),
		.PKT_TRANS_WRITE           (59),
		.PKT_TRANS_READ            (60),
		.OUT_NARROW_SIZE           (0),
		.IN_NARROW_SIZE            (1),
		.OUT_FIXED                 (0),
		.OUT_COMPLETE_WRAP         (0),
		.ST_DATA_W                 (113),
		.ST_CHANNEL_W              (8),
		.OUT_BYTE_CNT_H            (65),
		.OUT_BURSTWRAP_H           (76),
		.COMPRESSED_READ_SUPPORT   (1),
		.BYTEENABLE_SYNTHESIS      (1),
		.PIPE_INPUTS               (0),
		.NO_WRAP_SUPPORT           (0),
		.BURSTWRAP_CONST_MASK      (0),
		.BURSTWRAP_CONST_VALUE     (0)
	) burst_adapter_007 (
		.clk                   (pll_audio_outclk0_clk),                   //       cr0.clk
		.reset                 (rst_controller_003_reset_out_reset),      // cr0_reset.reset
		.sink0_valid           (cmd_xbar_mux_009_src_valid),              //     sink0.valid
		.sink0_data            (cmd_xbar_mux_009_src_data),               //          .data
		.sink0_channel         (cmd_xbar_mux_009_src_channel),            //          .channel
		.sink0_startofpacket   (cmd_xbar_mux_009_src_startofpacket),      //          .startofpacket
		.sink0_endofpacket     (cmd_xbar_mux_009_src_endofpacket),        //          .endofpacket
		.sink0_ready           (cmd_xbar_mux_009_src_ready),              //          .ready
		.source0_valid         (burst_adapter_007_source0_valid),         //   source0.valid
		.source0_data          (burst_adapter_007_source0_data),          //          .data
		.source0_channel       (burst_adapter_007_source0_channel),       //          .channel
		.source0_startofpacket (burst_adapter_007_source0_startofpacket), //          .startofpacket
		.source0_endofpacket   (burst_adapter_007_source0_endofpacket),   //          .endofpacket
		.source0_ready         (burst_adapter_007_source0_ready)          //          .ready
	);

	altera_merlin_burst_adapter #(
		.PKT_ADDR_H                (49),
		.PKT_ADDR_L                (18),
		.PKT_BEGIN_BURST           (83),
		.PKT_BYTE_CNT_H            (66),
		.PKT_BYTE_CNT_L            (56),
		.PKT_BYTEEN_H              (17),
		.PKT_BYTEEN_L              (16),
		.PKT_BURST_SIZE_H          (78),
		.PKT_BURST_SIZE_L          (76),
		.PKT_BURST_TYPE_H          (80),
		.PKT_BURST_TYPE_L          (79),
		.PKT_BURSTWRAP_H           (75),
		.PKT_BURSTWRAP_L           (67),
		.PKT_TRANS_COMPRESSED_READ (50),
		.PKT_TRANS_WRITE           (52),
		.PKT_TRANS_READ            (53),
		.OUT_NARROW_SIZE           (0),
		.IN_NARROW_SIZE            (1),
		.OUT_FIXED                 (0),
		.OUT_COMPLETE_WRAP         (0),
		.ST_DATA_W                 (108),
		.ST_CHANNEL_W              (3),
		.OUT_BYTE_CNT_H            (57),
		.OUT_BURSTWRAP_H           (75),
		.COMPRESSED_READ_SUPPORT   (1),
		.BYTEENABLE_SYNTHESIS      (1),
		.PIPE_INPUTS               (0),
		.NO_WRAP_SUPPORT           (0),
		.BURSTWRAP_CONST_MASK      (0),
		.BURSTWRAP_CONST_VALUE     (0)
	) burst_adapter_008 (
		.clk                   (pll_sdram_outclk1_clk),                      //       cr0.clk
		.reset                 (rst_controller_001_reset_out_reset),         // cr0_reset.reset
		.sink0_valid           (width_adapter_003_cmd_source_valid),         //     sink0.valid
		.sink0_data            (width_adapter_003_cmd_source_data),          //          .data
		.sink0_channel         (width_adapter_003_cmd_source_channel),       //          .channel
		.sink0_startofpacket   (width_adapter_003_cmd_source_startofpacket), //          .startofpacket
		.sink0_endofpacket     (width_adapter_003_cmd_source_endofpacket),   //          .endofpacket
		.sink0_ready           (width_adapter_003_cmd_source_ready),         //          .ready
		.source0_valid         (burst_adapter_008_source0_valid),            //   source0.valid
		.source0_data          (burst_adapter_008_source0_data),             //          .data
		.source0_channel       (burst_adapter_008_source0_channel),          //          .channel
		.source0_startofpacket (burst_adapter_008_source0_startofpacket),    //          .startofpacket
		.source0_endofpacket   (burst_adapter_008_source0_endofpacket),      //          .endofpacket
		.source0_ready         (burst_adapter_008_source0_ready)             //          .ready
	);

	altera_merlin_combined_width_adapter #(
		.IN_PKT_ADDR_H                 (67),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (81),
		.IN_PKT_BYTE_CNT_L             (74),
		.IN_PKT_TRANS_COMPRESSED_READ  (68),
		.IN_PKT_BURSTWRAP_H            (89),
		.IN_PKT_BURSTWRAP_L            (82),
		.IN_PKT_BURST_SIZE_H           (92),
		.IN_PKT_BURST_SIZE_L           (90),
		.IN_PKT_RESPONSE_STATUS_H      (114),
		.IN_PKT_RESPONSE_STATUS_L      (113),
		.IN_PKT_TRANS_EXCLUSIVE        (73),
		.IN_PKT_BURST_TYPE_H           (94),
		.IN_PKT_BURST_TYPE_L           (93),
		.IN_PKT_TRANS_POSTED           (69),
		.IN_ST_DATA_W                  (115),
		.OUT_PKT_ADDR_H                (103),
		.OUT_PKT_ADDR_L                (72),
		.OUT_PKT_DATA_H                (63),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (71),
		.OUT_PKT_BYTEEN_L              (64),
		.OUT_PKT_BYTE_CNT_H            (117),
		.OUT_PKT_BYTE_CNT_L            (110),
		.OUT_PKT_TRANS_COMPRESSED_READ (104),
		.OUT_PKT_TRANS_EXCLUSIVE       (109),
		.OUT_PKT_RESPONSE_STATUS_H     (150),
		.OUT_PKT_RESPONSE_STATUS_L     (149),
		.OUT_PKT_BURST_SIZE_H          (128),
		.OUT_PKT_BURST_SIZE_L          (126),
		.OUT_PKT_BURST_TYPE_H          (130),
		.OUT_PKT_BURST_TYPE_L          (129),
		.OUT_ST_DATA_W                 (151),
		.ST_CHANNEL_W                  (2),
		.MAX_OUTSTANDING_RESPONSES     (24)
	) width_adapter (
		.clk                   (clk_clk),                                //      clock.clk
		.reset                 (rst_controller_004_reset_out_reset),     //      reset.reset
		.cmd_in_valid          (cmd_xbar_demux_src0_valid),              //   cmd_sink.valid
		.cmd_in_channel        (cmd_xbar_demux_src0_channel),            //           .channel
		.cmd_in_data           (cmd_xbar_demux_src0_data),               //           .data
		.cmd_in_startofpacket  (cmd_xbar_demux_src0_startofpacket),      //           .startofpacket
		.cmd_in_endofpacket    (cmd_xbar_demux_src0_endofpacket),        //           .endofpacket
		.cmd_in_ready          (cmd_xbar_demux_src0_ready),              //           .ready
		.cmd_out_ready         (width_adapter_cmd_source_ready),         // cmd_source.ready
		.cmd_out_valid         (width_adapter_cmd_source_valid),         //           .valid
		.cmd_out_channel       (width_adapter_cmd_source_channel),       //           .channel
		.cmd_out_data          (width_adapter_cmd_source_data),          //           .data
		.cmd_out_startofpacket (width_adapter_cmd_source_startofpacket), //           .startofpacket
		.cmd_out_endofpacket   (width_adapter_cmd_source_endofpacket),   //           .endofpacket
		.rsp_in_ready          (id_router_src_ready),                    //   rsp_sink.ready
		.rsp_in_valid          (id_router_src_valid),                    //           .valid
		.rsp_in_channel        (id_router_src_channel),                  //           .channel
		.rsp_in_data           (id_router_src_data),                     //           .data
		.rsp_in_startofpacket  (id_router_src_startofpacket),            //           .startofpacket
		.rsp_in_endofpacket    (id_router_src_endofpacket),              //           .endofpacket
		.rsp_out_ready         (width_adapter_rsp_source_ready),         // rsp_source.ready
		.rsp_out_valid         (width_adapter_rsp_source_valid),         //           .valid
		.rsp_out_channel       (width_adapter_rsp_source_channel),       //           .channel
		.rsp_out_data          (width_adapter_rsp_source_data),          //           .data
		.rsp_out_startofpacket (width_adapter_rsp_source_startofpacket), //           .startofpacket
		.rsp_out_endofpacket   (width_adapter_rsp_source_endofpacket)    //           .endofpacket
	);

	altera_merlin_combined_width_adapter #(
		.IN_PKT_ADDR_H                 (67),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (81),
		.IN_PKT_BYTE_CNT_L             (74),
		.IN_PKT_TRANS_COMPRESSED_READ  (68),
		.IN_PKT_BURSTWRAP_H            (89),
		.IN_PKT_BURSTWRAP_L            (82),
		.IN_PKT_BURST_SIZE_H           (92),
		.IN_PKT_BURST_SIZE_L           (90),
		.IN_PKT_RESPONSE_STATUS_H      (114),
		.IN_PKT_RESPONSE_STATUS_L      (113),
		.IN_PKT_TRANS_EXCLUSIVE        (73),
		.IN_PKT_BURST_TYPE_H           (94),
		.IN_PKT_BURST_TYPE_L           (93),
		.IN_PKT_TRANS_POSTED           (69),
		.IN_ST_DATA_W                  (115),
		.OUT_PKT_ADDR_H                (103),
		.OUT_PKT_ADDR_L                (72),
		.OUT_PKT_DATA_H                (63),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (71),
		.OUT_PKT_BYTEEN_L              (64),
		.OUT_PKT_BYTE_CNT_H            (117),
		.OUT_PKT_BYTE_CNT_L            (110),
		.OUT_PKT_TRANS_COMPRESSED_READ (104),
		.OUT_PKT_TRANS_EXCLUSIVE       (109),
		.OUT_PKT_RESPONSE_STATUS_H     (150),
		.OUT_PKT_RESPONSE_STATUS_L     (149),
		.OUT_PKT_BURST_SIZE_H          (128),
		.OUT_PKT_BURST_SIZE_L          (126),
		.OUT_PKT_BURST_TYPE_H          (130),
		.OUT_PKT_BURST_TYPE_L          (129),
		.OUT_ST_DATA_W                 (151),
		.ST_CHANNEL_W                  (2),
		.MAX_OUTSTANDING_RESPONSES     (24)
	) width_adapter_001 (
		.clk                   (clk_clk),                                    //      clock.clk
		.reset                 (rst_controller_004_reset_out_reset),         //      reset.reset
		.cmd_in_valid          (cmd_xbar_demux_src1_valid),                  //   cmd_sink.valid
		.cmd_in_channel        (cmd_xbar_demux_src1_channel),                //           .channel
		.cmd_in_data           (cmd_xbar_demux_src1_data),                   //           .data
		.cmd_in_startofpacket  (cmd_xbar_demux_src1_startofpacket),          //           .startofpacket
		.cmd_in_endofpacket    (cmd_xbar_demux_src1_endofpacket),            //           .endofpacket
		.cmd_in_ready          (cmd_xbar_demux_src1_ready),                  //           .ready
		.cmd_out_ready         (width_adapter_001_cmd_source_ready),         // cmd_source.ready
		.cmd_out_valid         (width_adapter_001_cmd_source_valid),         //           .valid
		.cmd_out_channel       (width_adapter_001_cmd_source_channel),       //           .channel
		.cmd_out_data          (width_adapter_001_cmd_source_data),          //           .data
		.cmd_out_startofpacket (width_adapter_001_cmd_source_startofpacket), //           .startofpacket
		.cmd_out_endofpacket   (width_adapter_001_cmd_source_endofpacket),   //           .endofpacket
		.rsp_in_ready          (id_router_001_src_ready),                    //   rsp_sink.ready
		.rsp_in_valid          (id_router_001_src_valid),                    //           .valid
		.rsp_in_channel        (id_router_001_src_channel),                  //           .channel
		.rsp_in_data           (id_router_001_src_data),                     //           .data
		.rsp_in_startofpacket  (id_router_001_src_startofpacket),            //           .startofpacket
		.rsp_in_endofpacket    (id_router_001_src_endofpacket),              //           .endofpacket
		.rsp_out_ready         (width_adapter_001_rsp_source_ready),         // rsp_source.ready
		.rsp_out_valid         (width_adapter_001_rsp_source_valid),         //           .valid
		.rsp_out_channel       (width_adapter_001_rsp_source_channel),       //           .channel
		.rsp_out_data          (width_adapter_001_rsp_source_data),          //           .data
		.rsp_out_startofpacket (width_adapter_001_rsp_source_startofpacket), //           .startofpacket
		.rsp_out_endofpacket   (width_adapter_001_rsp_source_endofpacket)    //           .endofpacket
	);

	altera_merlin_combined_width_adapter #(
		.IN_PKT_ADDR_H                 (67),
		.IN_PKT_ADDR_L                 (36),
		.IN_PKT_DATA_H                 (31),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (35),
		.IN_PKT_BYTEEN_L               (32),
		.IN_PKT_BYTE_CNT_H             (84),
		.IN_PKT_BYTE_CNT_L             (74),
		.IN_PKT_TRANS_COMPRESSED_READ  (68),
		.IN_PKT_BURSTWRAP_H            (93),
		.IN_PKT_BURSTWRAP_L            (85),
		.IN_PKT_BURST_SIZE_H           (96),
		.IN_PKT_BURST_SIZE_L           (94),
		.IN_PKT_RESPONSE_STATUS_H      (125),
		.IN_PKT_RESPONSE_STATUS_L      (124),
		.IN_PKT_TRANS_EXCLUSIVE        (73),
		.IN_PKT_BURST_TYPE_H           (98),
		.IN_PKT_BURST_TYPE_L           (97),
		.IN_PKT_TRANS_POSTED           (69),
		.IN_ST_DATA_W                  (126),
		.OUT_PKT_ADDR_H                (175),
		.OUT_PKT_ADDR_L                (144),
		.OUT_PKT_DATA_H                (127),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (143),
		.OUT_PKT_BYTEEN_L              (128),
		.OUT_PKT_BYTE_CNT_H            (192),
		.OUT_PKT_BYTE_CNT_L            (182),
		.OUT_PKT_TRANS_COMPRESSED_READ (176),
		.OUT_PKT_TRANS_EXCLUSIVE       (181),
		.OUT_PKT_RESPONSE_STATUS_H     (233),
		.OUT_PKT_RESPONSE_STATUS_L     (232),
		.OUT_PKT_BURST_SIZE_H          (204),
		.OUT_PKT_BURST_SIZE_L          (202),
		.OUT_PKT_BURST_TYPE_H          (206),
		.OUT_PKT_BURST_TYPE_L          (205),
		.OUT_ST_DATA_W                 (234),
		.ST_CHANNEL_W                  (3),
		.MAX_OUTSTANDING_RESPONSES     (24)
	) width_adapter_002 (
		.clk                   (pll_sdram_outclk1_clk),                      //      clock.clk
		.reset                 (rst_controller_001_reset_out_reset),         //      reset.reset
		.cmd_in_valid          (addr_router_005_src_valid),                  //   cmd_sink.valid
		.cmd_in_channel        (addr_router_005_src_channel),                //           .channel
		.cmd_in_data           (addr_router_005_src_data),                   //           .data
		.cmd_in_startofpacket  (addr_router_005_src_startofpacket),          //           .startofpacket
		.cmd_in_endofpacket    (addr_router_005_src_endofpacket),            //           .endofpacket
		.cmd_in_ready          (addr_router_005_src_ready),                  //           .ready
		.cmd_out_ready         (width_adapter_002_cmd_source_ready),         // cmd_source.ready
		.cmd_out_valid         (width_adapter_002_cmd_source_valid),         //           .valid
		.cmd_out_channel       (width_adapter_002_cmd_source_channel),       //           .channel
		.cmd_out_data          (width_adapter_002_cmd_source_data),          //           .data
		.cmd_out_startofpacket (width_adapter_002_cmd_source_startofpacket), //           .startofpacket
		.cmd_out_endofpacket   (width_adapter_002_cmd_source_endofpacket),   //           .endofpacket
		.rsp_in_ready          (rsp_xbar_demux_010_src2_ready),              //   rsp_sink.ready
		.rsp_in_valid          (rsp_xbar_demux_010_src2_valid),              //           .valid
		.rsp_in_channel        (rsp_xbar_demux_010_src2_channel),            //           .channel
		.rsp_in_data           (rsp_xbar_demux_010_src2_data),               //           .data
		.rsp_in_startofpacket  (rsp_xbar_demux_010_src2_startofpacket),      //           .startofpacket
		.rsp_in_endofpacket    (rsp_xbar_demux_010_src2_endofpacket),        //           .endofpacket
		.rsp_out_ready         (width_adapter_002_rsp_source_ready),         // rsp_source.ready
		.rsp_out_valid         (width_adapter_002_rsp_source_valid),         //           .valid
		.rsp_out_channel       (width_adapter_002_rsp_source_channel),       //           .channel
		.rsp_out_data          (width_adapter_002_rsp_source_data),          //           .data
		.rsp_out_startofpacket (width_adapter_002_rsp_source_startofpacket), //           .startofpacket
		.rsp_out_endofpacket   (width_adapter_002_rsp_source_endofpacket)    //           .endofpacket
	);

	altera_merlin_combined_width_adapter #(
		.IN_PKT_ADDR_H                 (175),
		.IN_PKT_ADDR_L                 (144),
		.IN_PKT_DATA_H                 (127),
		.IN_PKT_DATA_L                 (0),
		.IN_PKT_BYTEEN_H               (143),
		.IN_PKT_BYTEEN_L               (128),
		.IN_PKT_BYTE_CNT_H             (192),
		.IN_PKT_BYTE_CNT_L             (182),
		.IN_PKT_TRANS_COMPRESSED_READ  (176),
		.IN_PKT_BURSTWRAP_H            (201),
		.IN_PKT_BURSTWRAP_L            (193),
		.IN_PKT_BURST_SIZE_H           (204),
		.IN_PKT_BURST_SIZE_L           (202),
		.IN_PKT_RESPONSE_STATUS_H      (233),
		.IN_PKT_RESPONSE_STATUS_L      (232),
		.IN_PKT_TRANS_EXCLUSIVE        (181),
		.IN_PKT_BURST_TYPE_H           (206),
		.IN_PKT_BURST_TYPE_L           (205),
		.IN_PKT_TRANS_POSTED           (177),
		.IN_ST_DATA_W                  (234),
		.OUT_PKT_ADDR_H                (49),
		.OUT_PKT_ADDR_L                (18),
		.OUT_PKT_DATA_H                (15),
		.OUT_PKT_DATA_L                (0),
		.OUT_PKT_BYTEEN_H              (17),
		.OUT_PKT_BYTEEN_L              (16),
		.OUT_PKT_BYTE_CNT_H            (66),
		.OUT_PKT_BYTE_CNT_L            (56),
		.OUT_PKT_TRANS_COMPRESSED_READ (50),
		.OUT_PKT_TRANS_EXCLUSIVE       (55),
		.OUT_PKT_RESPONSE_STATUS_H     (107),
		.OUT_PKT_RESPONSE_STATUS_L     (106),
		.OUT_PKT_BURST_SIZE_H          (78),
		.OUT_PKT_BURST_SIZE_L          (76),
		.OUT_PKT_BURST_TYPE_H          (80),
		.OUT_PKT_BURST_TYPE_L          (79),
		.OUT_ST_DATA_W                 (108),
		.ST_CHANNEL_W                  (3),
		.MAX_OUTSTANDING_RESPONSES     (24)
	) width_adapter_003 (
		.clk                   (pll_sdram_outclk1_clk),                      //      clock.clk
		.reset                 (rst_controller_001_reset_out_reset),         //      reset.reset
		.cmd_in_valid          (cmd_xbar_mux_010_src_valid),                 //   cmd_sink.valid
		.cmd_in_channel        (cmd_xbar_mux_010_src_channel),               //           .channel
		.cmd_in_data           (cmd_xbar_mux_010_src_data),                  //           .data
		.cmd_in_startofpacket  (cmd_xbar_mux_010_src_startofpacket),         //           .startofpacket
		.cmd_in_endofpacket    (cmd_xbar_mux_010_src_endofpacket),           //           .endofpacket
		.cmd_in_ready          (cmd_xbar_mux_010_src_ready),                 //           .ready
		.cmd_out_ready         (width_adapter_003_cmd_source_ready),         // cmd_source.ready
		.cmd_out_valid         (width_adapter_003_cmd_source_valid),         //           .valid
		.cmd_out_channel       (width_adapter_003_cmd_source_channel),       //           .channel
		.cmd_out_data          (width_adapter_003_cmd_source_data),          //           .data
		.cmd_out_startofpacket (width_adapter_003_cmd_source_startofpacket), //           .startofpacket
		.cmd_out_endofpacket   (width_adapter_003_cmd_source_endofpacket),   //           .endofpacket
		.rsp_in_ready          (id_router_010_src_ready),                    //   rsp_sink.ready
		.rsp_in_valid          (id_router_010_src_valid),                    //           .valid
		.rsp_in_channel        (id_router_010_src_channel),                  //           .channel
		.rsp_in_data           (id_router_010_src_data),                     //           .data
		.rsp_in_startofpacket  (id_router_010_src_startofpacket),            //           .startofpacket
		.rsp_in_endofpacket    (id_router_010_src_endofpacket),              //           .endofpacket
		.rsp_out_ready         (width_adapter_003_rsp_source_ready),         // rsp_source.ready
		.rsp_out_valid         (width_adapter_003_rsp_source_valid),         //           .valid
		.rsp_out_channel       (width_adapter_003_rsp_source_channel),       //           .channel
		.rsp_out_data          (width_adapter_003_rsp_source_data),          //           .data
		.rsp_out_startofpacket (width_adapter_003_rsp_source_startofpacket), //           .startofpacket
		.rsp_out_endofpacket   (width_adapter_003_rsp_source_endofpacket)    //           .endofpacket
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (1),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2),
		.RESET_REQUEST_PRESENT   (0)
	) rst_controller (
		.reset_in0  (~reset_reset_n),                 // reset_in0.reset
		.clk        (clk_clk),                        //       clk.clk
		.reset_out  (rst_controller_reset_out_reset), // reset_out.reset
		.reset_req  (),                               // (terminated)
		.reset_in1  (1'b0),                           // (terminated)
		.reset_in2  (1'b0),                           // (terminated)
		.reset_in3  (1'b0),                           // (terminated)
		.reset_in4  (1'b0),                           // (terminated)
		.reset_in5  (1'b0),                           // (terminated)
		.reset_in6  (1'b0),                           // (terminated)
		.reset_in7  (1'b0),                           // (terminated)
		.reset_in8  (1'b0),                           // (terminated)
		.reset_in9  (1'b0),                           // (terminated)
		.reset_in10 (1'b0),                           // (terminated)
		.reset_in11 (1'b0),                           // (terminated)
		.reset_in12 (1'b0),                           // (terminated)
		.reset_in13 (1'b0),                           // (terminated)
		.reset_in14 (1'b0),                           // (terminated)
		.reset_in15 (1'b0)                            // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (1),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2),
		.RESET_REQUEST_PRESENT   (0)
	) rst_controller_001 (
		.reset_in0  (~reset_reset_n),                     // reset_in0.reset
		.clk        (pll_sdram_outclk1_clk),              //       clk.clk
		.reset_out  (rst_controller_001_reset_out_reset), // reset_out.reset
		.reset_req  (),                                   // (terminated)
		.reset_in1  (1'b0),                               // (terminated)
		.reset_in2  (1'b0),                               // (terminated)
		.reset_in3  (1'b0),                               // (terminated)
		.reset_in4  (1'b0),                               // (terminated)
		.reset_in5  (1'b0),                               // (terminated)
		.reset_in6  (1'b0),                               // (terminated)
		.reset_in7  (1'b0),                               // (terminated)
		.reset_in8  (1'b0),                               // (terminated)
		.reset_in9  (1'b0),                               // (terminated)
		.reset_in10 (1'b0),                               // (terminated)
		.reset_in11 (1'b0),                               // (terminated)
		.reset_in12 (1'b0),                               // (terminated)
		.reset_in13 (1'b0),                               // (terminated)
		.reset_in14 (1'b0),                               // (terminated)
		.reset_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (1),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2),
		.RESET_REQUEST_PRESENT   (0)
	) rst_controller_002 (
		.reset_in0  (~reset_reset_n),                     // reset_in0.reset
		.clk        (pll_stream_outclk1_clk),             //       clk.clk
		.reset_out  (rst_controller_002_reset_out_reset), // reset_out.reset
		.reset_req  (),                                   // (terminated)
		.reset_in1  (1'b0),                               // (terminated)
		.reset_in2  (1'b0),                               // (terminated)
		.reset_in3  (1'b0),                               // (terminated)
		.reset_in4  (1'b0),                               // (terminated)
		.reset_in5  (1'b0),                               // (terminated)
		.reset_in6  (1'b0),                               // (terminated)
		.reset_in7  (1'b0),                               // (terminated)
		.reset_in8  (1'b0),                               // (terminated)
		.reset_in9  (1'b0),                               // (terminated)
		.reset_in10 (1'b0),                               // (terminated)
		.reset_in11 (1'b0),                               // (terminated)
		.reset_in12 (1'b0),                               // (terminated)
		.reset_in13 (1'b0),                               // (terminated)
		.reset_in14 (1'b0),                               // (terminated)
		.reset_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (1),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2),
		.RESET_REQUEST_PRESENT   (0)
	) rst_controller_003 (
		.reset_in0  (~reset_reset_n),                     // reset_in0.reset
		.clk        (pll_audio_outclk0_clk),              //       clk.clk
		.reset_out  (rst_controller_003_reset_out_reset), // reset_out.reset
		.reset_req  (),                                   // (terminated)
		.reset_in1  (1'b0),                               // (terminated)
		.reset_in2  (1'b0),                               // (terminated)
		.reset_in3  (1'b0),                               // (terminated)
		.reset_in4  (1'b0),                               // (terminated)
		.reset_in5  (1'b0),                               // (terminated)
		.reset_in6  (1'b0),                               // (terminated)
		.reset_in7  (1'b0),                               // (terminated)
		.reset_in8  (1'b0),                               // (terminated)
		.reset_in9  (1'b0),                               // (terminated)
		.reset_in10 (1'b0),                               // (terminated)
		.reset_in11 (1'b0),                               // (terminated)
		.reset_in12 (1'b0),                               // (terminated)
		.reset_in13 (1'b0),                               // (terminated)
		.reset_in14 (1'b0),                               // (terminated)
		.reset_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (1),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2),
		.RESET_REQUEST_PRESENT   (0)
	) rst_controller_004 (
		.reset_in0  (~hps_0_h2f_reset_reset_n),           // reset_in0.reset
		.clk        (clk_clk),                            //       clk.clk
		.reset_out  (rst_controller_004_reset_out_reset), // reset_out.reset
		.reset_req  (),                                   // (terminated)
		.reset_in1  (1'b0),                               // (terminated)
		.reset_in2  (1'b0),                               // (terminated)
		.reset_in3  (1'b0),                               // (terminated)
		.reset_in4  (1'b0),                               // (terminated)
		.reset_in5  (1'b0),                               // (terminated)
		.reset_in6  (1'b0),                               // (terminated)
		.reset_in7  (1'b0),                               // (terminated)
		.reset_in8  (1'b0),                               // (terminated)
		.reset_in9  (1'b0),                               // (terminated)
		.reset_in10 (1'b0),                               // (terminated)
		.reset_in11 (1'b0),                               // (terminated)
		.reset_in12 (1'b0),                               // (terminated)
		.reset_in13 (1'b0),                               // (terminated)
		.reset_in14 (1'b0),                               // (terminated)
		.reset_in15 (1'b0)                                // (terminated)
	);

	altera_reset_controller #(
		.NUM_RESET_INPUTS        (1),
		.OUTPUT_RESET_SYNC_EDGES ("deassert"),
		.SYNC_DEPTH              (2),
		.RESET_REQUEST_PRESENT   (0)
	) rst_controller_005 (
		.reset_in0  (~hps_0_h2f_reset_reset_n),           // reset_in0.reset
		.clk        (pll_sdram_outclk1_clk),              //       clk.clk
		.reset_out  (rst_controller_005_reset_out_reset), // reset_out.reset
		.reset_req  (),                                   // (terminated)
		.reset_in1  (1'b0),                               // (terminated)
		.reset_in2  (1'b0),                               // (terminated)
		.reset_in3  (1'b0),                               // (terminated)
		.reset_in4  (1'b0),                               // (terminated)
		.reset_in5  (1'b0),                               // (terminated)
		.reset_in6  (1'b0),                               // (terminated)
		.reset_in7  (1'b0),                               // (terminated)
		.reset_in8  (1'b0),                               // (terminated)
		.reset_in9  (1'b0),                               // (terminated)
		.reset_in10 (1'b0),                               // (terminated)
		.reset_in11 (1'b0),                               // (terminated)
		.reset_in12 (1'b0),                               // (terminated)
		.reset_in13 (1'b0),                               // (terminated)
		.reset_in14 (1'b0),                               // (terminated)
		.reset_in15 (1'b0)                                // (terminated)
	);

	soc_system_cmd_xbar_demux cmd_xbar_demux (
		.clk                (clk_clk),                           //        clk.clk
		.reset              (rst_controller_reset_out_reset),    //  clk_reset.reset
		.sink_ready         (limiter_cmd_src_ready),             //       sink.ready
		.sink_channel       (limiter_cmd_src_channel),           //           .channel
		.sink_data          (limiter_cmd_src_data),              //           .data
		.sink_startofpacket (limiter_cmd_src_startofpacket),     //           .startofpacket
		.sink_endofpacket   (limiter_cmd_src_endofpacket),       //           .endofpacket
		.sink_valid         (limiter_cmd_valid_data),            // sink_valid.data
		.src0_ready         (cmd_xbar_demux_src0_ready),         //       src0.ready
		.src0_valid         (cmd_xbar_demux_src0_valid),         //           .valid
		.src0_data          (cmd_xbar_demux_src0_data),          //           .data
		.src0_channel       (cmd_xbar_demux_src0_channel),       //           .channel
		.src0_startofpacket (cmd_xbar_demux_src0_startofpacket), //           .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_src0_endofpacket),   //           .endofpacket
		.src1_ready         (cmd_xbar_demux_src1_ready),         //       src1.ready
		.src1_valid         (cmd_xbar_demux_src1_valid),         //           .valid
		.src1_data          (cmd_xbar_demux_src1_data),          //           .data
		.src1_channel       (cmd_xbar_demux_src1_channel),       //           .channel
		.src1_startofpacket (cmd_xbar_demux_src1_startofpacket), //           .startofpacket
		.src1_endofpacket   (cmd_xbar_demux_src1_endofpacket)    //           .endofpacket
	);

	soc_system_rsp_xbar_demux rsp_xbar_demux (
		.clk                (clk_clk),                                //       clk.clk
		.reset              (rst_controller_004_reset_out_reset),     // clk_reset.reset
		.sink_ready         (width_adapter_rsp_source_ready),         //      sink.ready
		.sink_channel       (width_adapter_rsp_source_channel),       //          .channel
		.sink_data          (width_adapter_rsp_source_data),          //          .data
		.sink_startofpacket (width_adapter_rsp_source_startofpacket), //          .startofpacket
		.sink_endofpacket   (width_adapter_rsp_source_endofpacket),   //          .endofpacket
		.sink_valid         (width_adapter_rsp_source_valid),         //          .valid
		.src0_ready         (rsp_xbar_demux_src0_ready),              //      src0.ready
		.src0_valid         (rsp_xbar_demux_src0_valid),              //          .valid
		.src0_data          (rsp_xbar_demux_src0_data),               //          .data
		.src0_channel       (rsp_xbar_demux_src0_channel),            //          .channel
		.src0_startofpacket (rsp_xbar_demux_src0_startofpacket),      //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_src0_endofpacket)         //          .endofpacket
	);

	soc_system_rsp_xbar_demux rsp_xbar_demux_001 (
		.clk                (clk_clk),                                    //       clk.clk
		.reset              (rst_controller_004_reset_out_reset),         // clk_reset.reset
		.sink_ready         (width_adapter_001_rsp_source_ready),         //      sink.ready
		.sink_channel       (width_adapter_001_rsp_source_channel),       //          .channel
		.sink_data          (width_adapter_001_rsp_source_data),          //          .data
		.sink_startofpacket (width_adapter_001_rsp_source_startofpacket), //          .startofpacket
		.sink_endofpacket   (width_adapter_001_rsp_source_endofpacket),   //          .endofpacket
		.sink_valid         (width_adapter_001_rsp_source_valid),         //          .valid
		.src0_ready         (rsp_xbar_demux_001_src0_ready),              //      src0.ready
		.src0_valid         (rsp_xbar_demux_001_src0_valid),              //          .valid
		.src0_data          (rsp_xbar_demux_001_src0_data),               //          .data
		.src0_channel       (rsp_xbar_demux_001_src0_channel),            //          .channel
		.src0_startofpacket (rsp_xbar_demux_001_src0_startofpacket),      //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_001_src0_endofpacket)         //          .endofpacket
	);

	soc_system_rsp_xbar_mux rsp_xbar_mux (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (rsp_xbar_mux_src_ready),                //       src.ready
		.src_valid           (rsp_xbar_mux_src_valid),                //          .valid
		.src_data            (rsp_xbar_mux_src_data),                 //          .data
		.src_channel         (rsp_xbar_mux_src_channel),              //          .channel
		.src_startofpacket   (rsp_xbar_mux_src_startofpacket),        //          .startofpacket
		.src_endofpacket     (rsp_xbar_mux_src_endofpacket),          //          .endofpacket
		.sink0_ready         (rsp_xbar_demux_src0_ready),             //     sink0.ready
		.sink0_valid         (rsp_xbar_demux_src0_valid),             //          .valid
		.sink0_channel       (rsp_xbar_demux_src0_channel),           //          .channel
		.sink0_data          (rsp_xbar_demux_src0_data),              //          .data
		.sink0_startofpacket (rsp_xbar_demux_src0_startofpacket),     //          .startofpacket
		.sink0_endofpacket   (rsp_xbar_demux_src0_endofpacket),       //          .endofpacket
		.sink1_ready         (rsp_xbar_demux_001_src0_ready),         //     sink1.ready
		.sink1_valid         (rsp_xbar_demux_001_src0_valid),         //          .valid
		.sink1_channel       (rsp_xbar_demux_001_src0_channel),       //          .channel
		.sink1_data          (rsp_xbar_demux_001_src0_data),          //          .data
		.sink1_startofpacket (rsp_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (rsp_xbar_demux_001_src0_endofpacket)    //          .endofpacket
	);

	soc_system_cmd_xbar_demux_001 cmd_xbar_demux_001 (
		.clk                (clk_clk),                               //        clk.clk
		.reset              (rst_controller_004_reset_out_reset),    //  clk_reset.reset
		.sink_ready         (limiter_001_cmd_src_ready),             //       sink.ready
		.sink_channel       (limiter_001_cmd_src_channel),           //           .channel
		.sink_data          (limiter_001_cmd_src_data),              //           .data
		.sink_startofpacket (limiter_001_cmd_src_startofpacket),     //           .startofpacket
		.sink_endofpacket   (limiter_001_cmd_src_endofpacket),       //           .endofpacket
		.sink_valid         (limiter_001_cmd_valid_data),            // sink_valid.data
		.src0_ready         (cmd_xbar_demux_001_src0_ready),         //       src0.ready
		.src0_valid         (cmd_xbar_demux_001_src0_valid),         //           .valid
		.src0_data          (cmd_xbar_demux_001_src0_data),          //           .data
		.src0_channel       (cmd_xbar_demux_001_src0_channel),       //           .channel
		.src0_startofpacket (cmd_xbar_demux_001_src0_startofpacket), //           .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_001_src0_endofpacket),   //           .endofpacket
		.src1_ready         (cmd_xbar_demux_001_src1_ready),         //       src1.ready
		.src1_valid         (cmd_xbar_demux_001_src1_valid),         //           .valid
		.src1_data          (cmd_xbar_demux_001_src1_data),          //           .data
		.src1_channel       (cmd_xbar_demux_001_src1_channel),       //           .channel
		.src1_startofpacket (cmd_xbar_demux_001_src1_startofpacket), //           .startofpacket
		.src1_endofpacket   (cmd_xbar_demux_001_src1_endofpacket),   //           .endofpacket
		.src2_ready         (cmd_xbar_demux_001_src2_ready),         //       src2.ready
		.src2_valid         (cmd_xbar_demux_001_src2_valid),         //           .valid
		.src2_data          (cmd_xbar_demux_001_src2_data),          //           .data
		.src2_channel       (cmd_xbar_demux_001_src2_channel),       //           .channel
		.src2_startofpacket (cmd_xbar_demux_001_src2_startofpacket), //           .startofpacket
		.src2_endofpacket   (cmd_xbar_demux_001_src2_endofpacket),   //           .endofpacket
		.src3_ready         (cmd_xbar_demux_001_src3_ready),         //       src3.ready
		.src3_valid         (cmd_xbar_demux_001_src3_valid),         //           .valid
		.src3_data          (cmd_xbar_demux_001_src3_data),          //           .data
		.src3_channel       (cmd_xbar_demux_001_src3_channel),       //           .channel
		.src3_startofpacket (cmd_xbar_demux_001_src3_startofpacket), //           .startofpacket
		.src3_endofpacket   (cmd_xbar_demux_001_src3_endofpacket),   //           .endofpacket
		.src4_ready         (cmd_xbar_demux_001_src4_ready),         //       src4.ready
		.src4_valid         (cmd_xbar_demux_001_src4_valid),         //           .valid
		.src4_data          (cmd_xbar_demux_001_src4_data),          //           .data
		.src4_channel       (cmd_xbar_demux_001_src4_channel),       //           .channel
		.src4_startofpacket (cmd_xbar_demux_001_src4_startofpacket), //           .startofpacket
		.src4_endofpacket   (cmd_xbar_demux_001_src4_endofpacket),   //           .endofpacket
		.src5_ready         (cmd_xbar_demux_001_src5_ready),         //       src5.ready
		.src5_valid         (cmd_xbar_demux_001_src5_valid),         //           .valid
		.src5_data          (cmd_xbar_demux_001_src5_data),          //           .data
		.src5_channel       (cmd_xbar_demux_001_src5_channel),       //           .channel
		.src5_startofpacket (cmd_xbar_demux_001_src5_startofpacket), //           .startofpacket
		.src5_endofpacket   (cmd_xbar_demux_001_src5_endofpacket),   //           .endofpacket
		.src6_ready         (cmd_xbar_demux_001_src6_ready),         //       src6.ready
		.src6_valid         (cmd_xbar_demux_001_src6_valid),         //           .valid
		.src6_data          (cmd_xbar_demux_001_src6_data),          //           .data
		.src6_channel       (cmd_xbar_demux_001_src6_channel),       //           .channel
		.src6_startofpacket (cmd_xbar_demux_001_src6_startofpacket), //           .startofpacket
		.src6_endofpacket   (cmd_xbar_demux_001_src6_endofpacket),   //           .endofpacket
		.src7_ready         (cmd_xbar_demux_001_src7_ready),         //       src7.ready
		.src7_valid         (cmd_xbar_demux_001_src7_valid),         //           .valid
		.src7_data          (cmd_xbar_demux_001_src7_data),          //           .data
		.src7_channel       (cmd_xbar_demux_001_src7_channel),       //           .channel
		.src7_startofpacket (cmd_xbar_demux_001_src7_startofpacket), //           .startofpacket
		.src7_endofpacket   (cmd_xbar_demux_001_src7_endofpacket)    //           .endofpacket
	);

	soc_system_cmd_xbar_demux_001 cmd_xbar_demux_002 (
		.clk                (clk_clk),                               //        clk.clk
		.reset              (rst_controller_004_reset_out_reset),    //  clk_reset.reset
		.sink_ready         (limiter_002_cmd_src_ready),             //       sink.ready
		.sink_channel       (limiter_002_cmd_src_channel),           //           .channel
		.sink_data          (limiter_002_cmd_src_data),              //           .data
		.sink_startofpacket (limiter_002_cmd_src_startofpacket),     //           .startofpacket
		.sink_endofpacket   (limiter_002_cmd_src_endofpacket),       //           .endofpacket
		.sink_valid         (limiter_002_cmd_valid_data),            // sink_valid.data
		.src0_ready         (cmd_xbar_demux_002_src0_ready),         //       src0.ready
		.src0_valid         (cmd_xbar_demux_002_src0_valid),         //           .valid
		.src0_data          (cmd_xbar_demux_002_src0_data),          //           .data
		.src0_channel       (cmd_xbar_demux_002_src0_channel),       //           .channel
		.src0_startofpacket (cmd_xbar_demux_002_src0_startofpacket), //           .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_002_src0_endofpacket),   //           .endofpacket
		.src1_ready         (cmd_xbar_demux_002_src1_ready),         //       src1.ready
		.src1_valid         (cmd_xbar_demux_002_src1_valid),         //           .valid
		.src1_data          (cmd_xbar_demux_002_src1_data),          //           .data
		.src1_channel       (cmd_xbar_demux_002_src1_channel),       //           .channel
		.src1_startofpacket (cmd_xbar_demux_002_src1_startofpacket), //           .startofpacket
		.src1_endofpacket   (cmd_xbar_demux_002_src1_endofpacket),   //           .endofpacket
		.src2_ready         (cmd_xbar_demux_002_src2_ready),         //       src2.ready
		.src2_valid         (cmd_xbar_demux_002_src2_valid),         //           .valid
		.src2_data          (cmd_xbar_demux_002_src2_data),          //           .data
		.src2_channel       (cmd_xbar_demux_002_src2_channel),       //           .channel
		.src2_startofpacket (cmd_xbar_demux_002_src2_startofpacket), //           .startofpacket
		.src2_endofpacket   (cmd_xbar_demux_002_src2_endofpacket),   //           .endofpacket
		.src3_ready         (cmd_xbar_demux_002_src3_ready),         //       src3.ready
		.src3_valid         (cmd_xbar_demux_002_src3_valid),         //           .valid
		.src3_data          (cmd_xbar_demux_002_src3_data),          //           .data
		.src3_channel       (cmd_xbar_demux_002_src3_channel),       //           .channel
		.src3_startofpacket (cmd_xbar_demux_002_src3_startofpacket), //           .startofpacket
		.src3_endofpacket   (cmd_xbar_demux_002_src3_endofpacket),   //           .endofpacket
		.src4_ready         (cmd_xbar_demux_002_src4_ready),         //       src4.ready
		.src4_valid         (cmd_xbar_demux_002_src4_valid),         //           .valid
		.src4_data          (cmd_xbar_demux_002_src4_data),          //           .data
		.src4_channel       (cmd_xbar_demux_002_src4_channel),       //           .channel
		.src4_startofpacket (cmd_xbar_demux_002_src4_startofpacket), //           .startofpacket
		.src4_endofpacket   (cmd_xbar_demux_002_src4_endofpacket),   //           .endofpacket
		.src5_ready         (cmd_xbar_demux_002_src5_ready),         //       src5.ready
		.src5_valid         (cmd_xbar_demux_002_src5_valid),         //           .valid
		.src5_data          (cmd_xbar_demux_002_src5_data),          //           .data
		.src5_channel       (cmd_xbar_demux_002_src5_channel),       //           .channel
		.src5_startofpacket (cmd_xbar_demux_002_src5_startofpacket), //           .startofpacket
		.src5_endofpacket   (cmd_xbar_demux_002_src5_endofpacket),   //           .endofpacket
		.src6_ready         (cmd_xbar_demux_002_src6_ready),         //       src6.ready
		.src6_valid         (cmd_xbar_demux_002_src6_valid),         //           .valid
		.src6_data          (cmd_xbar_demux_002_src6_data),          //           .data
		.src6_channel       (cmd_xbar_demux_002_src6_channel),       //           .channel
		.src6_startofpacket (cmd_xbar_demux_002_src6_startofpacket), //           .startofpacket
		.src6_endofpacket   (cmd_xbar_demux_002_src6_endofpacket),   //           .endofpacket
		.src7_ready         (cmd_xbar_demux_002_src7_ready),         //       src7.ready
		.src7_valid         (cmd_xbar_demux_002_src7_valid),         //           .valid
		.src7_data          (cmd_xbar_demux_002_src7_data),          //           .data
		.src7_channel       (cmd_xbar_demux_002_src7_channel),       //           .channel
		.src7_startofpacket (cmd_xbar_demux_002_src7_startofpacket), //           .startofpacket
		.src7_endofpacket   (cmd_xbar_demux_002_src7_endofpacket)    //           .endofpacket
	);

	soc_system_cmd_xbar_mux_002 cmd_xbar_mux_002 (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_002_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_002_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_002_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_002_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_002_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_002_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_001_src0_ready),         //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_001_src0_valid),         //          .valid
		.sink0_channel       (cmd_xbar_demux_001_src0_channel),       //          .channel
		.sink0_data          (cmd_xbar_demux_001_src0_data),          //          .data
		.sink0_startofpacket (cmd_xbar_demux_001_src0_startofpacket), //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_001_src0_endofpacket),   //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_002_src0_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_002_src0_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_002_src0_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_002_src0_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_002_src0_endofpacket)    //          .endofpacket
	);

	soc_system_cmd_xbar_mux_002 cmd_xbar_mux_003 (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_003_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_003_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_003_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_003_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_003_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_003_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_001_src1_ready),         //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_001_src1_valid),         //          .valid
		.sink0_channel       (cmd_xbar_demux_001_src1_channel),       //          .channel
		.sink0_data          (cmd_xbar_demux_001_src1_data),          //          .data
		.sink0_startofpacket (cmd_xbar_demux_001_src1_startofpacket), //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_001_src1_endofpacket),   //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_002_src1_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_002_src1_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_002_src1_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_002_src1_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_002_src1_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_002_src1_endofpacket)    //          .endofpacket
	);

	soc_system_cmd_xbar_mux_002 cmd_xbar_mux_004 (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_004_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_004_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_004_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_004_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_004_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_004_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_001_src2_ready),         //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_001_src2_valid),         //          .valid
		.sink0_channel       (cmd_xbar_demux_001_src2_channel),       //          .channel
		.sink0_data          (cmd_xbar_demux_001_src2_data),          //          .data
		.sink0_startofpacket (cmd_xbar_demux_001_src2_startofpacket), //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_001_src2_endofpacket),   //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_002_src2_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_002_src2_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_002_src2_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_002_src2_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_002_src2_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_002_src2_endofpacket)    //          .endofpacket
	);

	soc_system_cmd_xbar_mux_002 cmd_xbar_mux_005 (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_005_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_005_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_005_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_005_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_005_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_005_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_001_src3_ready),         //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_001_src3_valid),         //          .valid
		.sink0_channel       (cmd_xbar_demux_001_src3_channel),       //          .channel
		.sink0_data          (cmd_xbar_demux_001_src3_data),          //          .data
		.sink0_startofpacket (cmd_xbar_demux_001_src3_startofpacket), //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_001_src3_endofpacket),   //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_002_src3_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_002_src3_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_002_src3_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_002_src3_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_002_src3_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_002_src3_endofpacket)    //          .endofpacket
	);

	soc_system_cmd_xbar_mux_002 cmd_xbar_mux_006 (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_reset_out_reset),        // clk_reset.reset
		.src_ready           (cmd_xbar_mux_006_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_006_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_006_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_006_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_006_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_006_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_001_src4_ready),         //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_001_src4_valid),         //          .valid
		.sink0_channel       (cmd_xbar_demux_001_src4_channel),       //          .channel
		.sink0_data          (cmd_xbar_demux_001_src4_data),          //          .data
		.sink0_startofpacket (cmd_xbar_demux_001_src4_startofpacket), //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_001_src4_endofpacket),   //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_002_src4_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_002_src4_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_002_src4_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_002_src4_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_002_src4_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_002_src4_endofpacket)    //          .endofpacket
	);

	soc_system_cmd_xbar_mux_002 cmd_xbar_mux_007 (
		.clk                 (pll_stream_outclk1_clk),             //       clk.clk
		.reset               (rst_controller_002_reset_out_reset), // clk_reset.reset
		.src_ready           (cmd_xbar_mux_007_src_ready),         //       src.ready
		.src_valid           (cmd_xbar_mux_007_src_valid),         //          .valid
		.src_data            (cmd_xbar_mux_007_src_data),          //          .data
		.src_channel         (cmd_xbar_mux_007_src_channel),       //          .channel
		.src_startofpacket   (cmd_xbar_mux_007_src_startofpacket), //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_007_src_endofpacket),   //          .endofpacket
		.sink0_ready         (crosser_out_ready),                  //     sink0.ready
		.sink0_valid         (crosser_out_valid),                  //          .valid
		.sink0_channel       (crosser_out_channel),                //          .channel
		.sink0_data          (crosser_out_data),                   //          .data
		.sink0_startofpacket (crosser_out_startofpacket),          //          .startofpacket
		.sink0_endofpacket   (crosser_out_endofpacket),            //          .endofpacket
		.sink1_ready         (crosser_003_out_ready),              //     sink1.ready
		.sink1_valid         (crosser_003_out_valid),              //          .valid
		.sink1_channel       (crosser_003_out_channel),            //          .channel
		.sink1_data          (crosser_003_out_data),               //          .data
		.sink1_startofpacket (crosser_003_out_startofpacket),      //          .startofpacket
		.sink1_endofpacket   (crosser_003_out_endofpacket)         //          .endofpacket
	);

	soc_system_cmd_xbar_mux_002 cmd_xbar_mux_008 (
		.clk                 (pll_stream_outclk1_clk),             //       clk.clk
		.reset               (rst_controller_002_reset_out_reset), // clk_reset.reset
		.src_ready           (cmd_xbar_mux_008_src_ready),         //       src.ready
		.src_valid           (cmd_xbar_mux_008_src_valid),         //          .valid
		.src_data            (cmd_xbar_mux_008_src_data),          //          .data
		.src_channel         (cmd_xbar_mux_008_src_channel),       //          .channel
		.src_startofpacket   (cmd_xbar_mux_008_src_startofpacket), //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_008_src_endofpacket),   //          .endofpacket
		.sink0_ready         (crosser_001_out_ready),              //     sink0.ready
		.sink0_valid         (crosser_001_out_valid),              //          .valid
		.sink0_channel       (crosser_001_out_channel),            //          .channel
		.sink0_data          (crosser_001_out_data),               //          .data
		.sink0_startofpacket (crosser_001_out_startofpacket),      //          .startofpacket
		.sink0_endofpacket   (crosser_001_out_endofpacket),        //          .endofpacket
		.sink1_ready         (crosser_004_out_ready),              //     sink1.ready
		.sink1_valid         (crosser_004_out_valid),              //          .valid
		.sink1_channel       (crosser_004_out_channel),            //          .channel
		.sink1_data          (crosser_004_out_data),               //          .data
		.sink1_startofpacket (crosser_004_out_startofpacket),      //          .startofpacket
		.sink1_endofpacket   (crosser_004_out_endofpacket)         //          .endofpacket
	);

	soc_system_cmd_xbar_mux_002 cmd_xbar_mux_009 (
		.clk                 (pll_audio_outclk0_clk),              //       clk.clk
		.reset               (rst_controller_003_reset_out_reset), // clk_reset.reset
		.src_ready           (cmd_xbar_mux_009_src_ready),         //       src.ready
		.src_valid           (cmd_xbar_mux_009_src_valid),         //          .valid
		.src_data            (cmd_xbar_mux_009_src_data),          //          .data
		.src_channel         (cmd_xbar_mux_009_src_channel),       //          .channel
		.src_startofpacket   (cmd_xbar_mux_009_src_startofpacket), //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_009_src_endofpacket),   //          .endofpacket
		.sink0_ready         (crosser_002_out_ready),              //     sink0.ready
		.sink0_valid         (crosser_002_out_valid),              //          .valid
		.sink0_channel       (crosser_002_out_channel),            //          .channel
		.sink0_data          (crosser_002_out_data),               //          .data
		.sink0_startofpacket (crosser_002_out_startofpacket),      //          .startofpacket
		.sink0_endofpacket   (crosser_002_out_endofpacket),        //          .endofpacket
		.sink1_ready         (crosser_005_out_ready),              //     sink1.ready
		.sink1_valid         (crosser_005_out_valid),              //          .valid
		.sink1_channel       (crosser_005_out_channel),            //          .channel
		.sink1_data          (crosser_005_out_data),               //          .data
		.sink1_startofpacket (crosser_005_out_startofpacket),      //          .startofpacket
		.sink1_endofpacket   (crosser_005_out_endofpacket)         //          .endofpacket
	);

	soc_system_rsp_xbar_demux_002 rsp_xbar_demux_002 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_002_src_ready),               //      sink.ready
		.sink_channel       (id_router_002_src_channel),             //          .channel
		.sink_data          (id_router_002_src_data),                //          .data
		.sink_startofpacket (id_router_002_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_002_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_002_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_002_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_002_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_002_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_002_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_002_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_002_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_002_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_002_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_002_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_002_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_002_src1_endofpacket)    //          .endofpacket
	);

	soc_system_rsp_xbar_demux_002 rsp_xbar_demux_003 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_003_src_ready),               //      sink.ready
		.sink_channel       (id_router_003_src_channel),             //          .channel
		.sink_data          (id_router_003_src_data),                //          .data
		.sink_startofpacket (id_router_003_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_003_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_003_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_003_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_003_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_003_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_003_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_003_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_003_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_003_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_003_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_003_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_003_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_003_src1_endofpacket)    //          .endofpacket
	);

	soc_system_rsp_xbar_demux_002 rsp_xbar_demux_004 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_004_src_ready),               //      sink.ready
		.sink_channel       (id_router_004_src_channel),             //          .channel
		.sink_data          (id_router_004_src_data),                //          .data
		.sink_startofpacket (id_router_004_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_004_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_004_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_004_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_004_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_004_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_004_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_004_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_004_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_004_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_004_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_004_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_004_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_004_src1_endofpacket)    //          .endofpacket
	);

	soc_system_rsp_xbar_demux_002 rsp_xbar_demux_005 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_005_src_ready),               //      sink.ready
		.sink_channel       (id_router_005_src_channel),             //          .channel
		.sink_data          (id_router_005_src_data),                //          .data
		.sink_startofpacket (id_router_005_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_005_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_005_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_005_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_005_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_005_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_005_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_005_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_005_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_005_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_005_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_005_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_005_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_005_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_005_src1_endofpacket)    //          .endofpacket
	);

	soc_system_rsp_xbar_demux_002 rsp_xbar_demux_006 (
		.clk                (clk_clk),                               //       clk.clk
		.reset              (rst_controller_reset_out_reset),        // clk_reset.reset
		.sink_ready         (id_router_006_src_ready),               //      sink.ready
		.sink_channel       (id_router_006_src_channel),             //          .channel
		.sink_data          (id_router_006_src_data),                //          .data
		.sink_startofpacket (id_router_006_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_006_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_006_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_006_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_006_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_006_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_006_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_006_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_006_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_006_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_006_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_006_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_006_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_006_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_006_src1_endofpacket)    //          .endofpacket
	);

	soc_system_rsp_xbar_demux_002 rsp_xbar_demux_007 (
		.clk                (pll_stream_outclk1_clk),                //       clk.clk
		.reset              (rst_controller_002_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_007_src_ready),               //      sink.ready
		.sink_channel       (id_router_007_src_channel),             //          .channel
		.sink_data          (id_router_007_src_data),                //          .data
		.sink_startofpacket (id_router_007_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_007_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_007_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_007_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_007_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_007_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_007_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_007_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_007_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_007_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_007_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_007_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_007_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_007_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_007_src1_endofpacket)    //          .endofpacket
	);

	soc_system_rsp_xbar_demux_002 rsp_xbar_demux_008 (
		.clk                (pll_stream_outclk1_clk),                //       clk.clk
		.reset              (rst_controller_002_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_008_src_ready),               //      sink.ready
		.sink_channel       (id_router_008_src_channel),             //          .channel
		.sink_data          (id_router_008_src_data),                //          .data
		.sink_startofpacket (id_router_008_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_008_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_008_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_008_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_008_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_008_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_008_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_008_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_008_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_008_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_008_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_008_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_008_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_008_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_008_src1_endofpacket)    //          .endofpacket
	);

	soc_system_rsp_xbar_demux_002 rsp_xbar_demux_009 (
		.clk                (pll_audio_outclk0_clk),                 //       clk.clk
		.reset              (rst_controller_003_reset_out_reset),    // clk_reset.reset
		.sink_ready         (id_router_009_src_ready),               //      sink.ready
		.sink_channel       (id_router_009_src_channel),             //          .channel
		.sink_data          (id_router_009_src_data),                //          .data
		.sink_startofpacket (id_router_009_src_startofpacket),       //          .startofpacket
		.sink_endofpacket   (id_router_009_src_endofpacket),         //          .endofpacket
		.sink_valid         (id_router_009_src_valid),               //          .valid
		.src0_ready         (rsp_xbar_demux_009_src0_ready),         //      src0.ready
		.src0_valid         (rsp_xbar_demux_009_src0_valid),         //          .valid
		.src0_data          (rsp_xbar_demux_009_src0_data),          //          .data
		.src0_channel       (rsp_xbar_demux_009_src0_channel),       //          .channel
		.src0_startofpacket (rsp_xbar_demux_009_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_009_src0_endofpacket),   //          .endofpacket
		.src1_ready         (rsp_xbar_demux_009_src1_ready),         //      src1.ready
		.src1_valid         (rsp_xbar_demux_009_src1_valid),         //          .valid
		.src1_data          (rsp_xbar_demux_009_src1_data),          //          .data
		.src1_channel       (rsp_xbar_demux_009_src1_channel),       //          .channel
		.src1_startofpacket (rsp_xbar_demux_009_src1_startofpacket), //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_009_src1_endofpacket)    //          .endofpacket
	);

	soc_system_rsp_xbar_mux_001 rsp_xbar_mux_001 (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_004_reset_out_reset),    // clk_reset.reset
		.src_ready           (rsp_xbar_mux_001_src_ready),            //       src.ready
		.src_valid           (rsp_xbar_mux_001_src_valid),            //          .valid
		.src_data            (rsp_xbar_mux_001_src_data),             //          .data
		.src_channel         (rsp_xbar_mux_001_src_channel),          //          .channel
		.src_startofpacket   (rsp_xbar_mux_001_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (rsp_xbar_mux_001_src_endofpacket),      //          .endofpacket
		.sink0_ready         (rsp_xbar_demux_002_src0_ready),         //     sink0.ready
		.sink0_valid         (rsp_xbar_demux_002_src0_valid),         //          .valid
		.sink0_channel       (rsp_xbar_demux_002_src0_channel),       //          .channel
		.sink0_data          (rsp_xbar_demux_002_src0_data),          //          .data
		.sink0_startofpacket (rsp_xbar_demux_002_src0_startofpacket), //          .startofpacket
		.sink0_endofpacket   (rsp_xbar_demux_002_src0_endofpacket),   //          .endofpacket
		.sink1_ready         (rsp_xbar_demux_003_src0_ready),         //     sink1.ready
		.sink1_valid         (rsp_xbar_demux_003_src0_valid),         //          .valid
		.sink1_channel       (rsp_xbar_demux_003_src0_channel),       //          .channel
		.sink1_data          (rsp_xbar_demux_003_src0_data),          //          .data
		.sink1_startofpacket (rsp_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (rsp_xbar_demux_003_src0_endofpacket),   //          .endofpacket
		.sink2_ready         (rsp_xbar_demux_004_src0_ready),         //     sink2.ready
		.sink2_valid         (rsp_xbar_demux_004_src0_valid),         //          .valid
		.sink2_channel       (rsp_xbar_demux_004_src0_channel),       //          .channel
		.sink2_data          (rsp_xbar_demux_004_src0_data),          //          .data
		.sink2_startofpacket (rsp_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.sink2_endofpacket   (rsp_xbar_demux_004_src0_endofpacket),   //          .endofpacket
		.sink3_ready         (rsp_xbar_demux_005_src0_ready),         //     sink3.ready
		.sink3_valid         (rsp_xbar_demux_005_src0_valid),         //          .valid
		.sink3_channel       (rsp_xbar_demux_005_src0_channel),       //          .channel
		.sink3_data          (rsp_xbar_demux_005_src0_data),          //          .data
		.sink3_startofpacket (rsp_xbar_demux_005_src0_startofpacket), //          .startofpacket
		.sink3_endofpacket   (rsp_xbar_demux_005_src0_endofpacket),   //          .endofpacket
		.sink4_ready         (rsp_xbar_demux_006_src0_ready),         //     sink4.ready
		.sink4_valid         (rsp_xbar_demux_006_src0_valid),         //          .valid
		.sink4_channel       (rsp_xbar_demux_006_src0_channel),       //          .channel
		.sink4_data          (rsp_xbar_demux_006_src0_data),          //          .data
		.sink4_startofpacket (rsp_xbar_demux_006_src0_startofpacket), //          .startofpacket
		.sink4_endofpacket   (rsp_xbar_demux_006_src0_endofpacket),   //          .endofpacket
		.sink5_ready         (crosser_006_out_ready),                 //     sink5.ready
		.sink5_valid         (crosser_006_out_valid),                 //          .valid
		.sink5_channel       (crosser_006_out_channel),               //          .channel
		.sink5_data          (crosser_006_out_data),                  //          .data
		.sink5_startofpacket (crosser_006_out_startofpacket),         //          .startofpacket
		.sink5_endofpacket   (crosser_006_out_endofpacket),           //          .endofpacket
		.sink6_ready         (crosser_008_out_ready),                 //     sink6.ready
		.sink6_valid         (crosser_008_out_valid),                 //          .valid
		.sink6_channel       (crosser_008_out_channel),               //          .channel
		.sink6_data          (crosser_008_out_data),                  //          .data
		.sink6_startofpacket (crosser_008_out_startofpacket),         //          .startofpacket
		.sink6_endofpacket   (crosser_008_out_endofpacket),           //          .endofpacket
		.sink7_ready         (crosser_010_out_ready),                 //     sink7.ready
		.sink7_valid         (crosser_010_out_valid),                 //          .valid
		.sink7_channel       (crosser_010_out_channel),               //          .channel
		.sink7_data          (crosser_010_out_data),                  //          .data
		.sink7_startofpacket (crosser_010_out_startofpacket),         //          .startofpacket
		.sink7_endofpacket   (crosser_010_out_endofpacket)            //          .endofpacket
	);

	soc_system_rsp_xbar_mux_001 rsp_xbar_mux_002 (
		.clk                 (clk_clk),                               //       clk.clk
		.reset               (rst_controller_004_reset_out_reset),    // clk_reset.reset
		.src_ready           (rsp_xbar_mux_002_src_ready),            //       src.ready
		.src_valid           (rsp_xbar_mux_002_src_valid),            //          .valid
		.src_data            (rsp_xbar_mux_002_src_data),             //          .data
		.src_channel         (rsp_xbar_mux_002_src_channel),          //          .channel
		.src_startofpacket   (rsp_xbar_mux_002_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (rsp_xbar_mux_002_src_endofpacket),      //          .endofpacket
		.sink0_ready         (rsp_xbar_demux_002_src1_ready),         //     sink0.ready
		.sink0_valid         (rsp_xbar_demux_002_src1_valid),         //          .valid
		.sink0_channel       (rsp_xbar_demux_002_src1_channel),       //          .channel
		.sink0_data          (rsp_xbar_demux_002_src1_data),          //          .data
		.sink0_startofpacket (rsp_xbar_demux_002_src1_startofpacket), //          .startofpacket
		.sink0_endofpacket   (rsp_xbar_demux_002_src1_endofpacket),   //          .endofpacket
		.sink1_ready         (rsp_xbar_demux_003_src1_ready),         //     sink1.ready
		.sink1_valid         (rsp_xbar_demux_003_src1_valid),         //          .valid
		.sink1_channel       (rsp_xbar_demux_003_src1_channel),       //          .channel
		.sink1_data          (rsp_xbar_demux_003_src1_data),          //          .data
		.sink1_startofpacket (rsp_xbar_demux_003_src1_startofpacket), //          .startofpacket
		.sink1_endofpacket   (rsp_xbar_demux_003_src1_endofpacket),   //          .endofpacket
		.sink2_ready         (rsp_xbar_demux_004_src1_ready),         //     sink2.ready
		.sink2_valid         (rsp_xbar_demux_004_src1_valid),         //          .valid
		.sink2_channel       (rsp_xbar_demux_004_src1_channel),       //          .channel
		.sink2_data          (rsp_xbar_demux_004_src1_data),          //          .data
		.sink2_startofpacket (rsp_xbar_demux_004_src1_startofpacket), //          .startofpacket
		.sink2_endofpacket   (rsp_xbar_demux_004_src1_endofpacket),   //          .endofpacket
		.sink3_ready         (rsp_xbar_demux_005_src1_ready),         //     sink3.ready
		.sink3_valid         (rsp_xbar_demux_005_src1_valid),         //          .valid
		.sink3_channel       (rsp_xbar_demux_005_src1_channel),       //          .channel
		.sink3_data          (rsp_xbar_demux_005_src1_data),          //          .data
		.sink3_startofpacket (rsp_xbar_demux_005_src1_startofpacket), //          .startofpacket
		.sink3_endofpacket   (rsp_xbar_demux_005_src1_endofpacket),   //          .endofpacket
		.sink4_ready         (rsp_xbar_demux_006_src1_ready),         //     sink4.ready
		.sink4_valid         (rsp_xbar_demux_006_src1_valid),         //          .valid
		.sink4_channel       (rsp_xbar_demux_006_src1_channel),       //          .channel
		.sink4_data          (rsp_xbar_demux_006_src1_data),          //          .data
		.sink4_startofpacket (rsp_xbar_demux_006_src1_startofpacket), //          .startofpacket
		.sink4_endofpacket   (rsp_xbar_demux_006_src1_endofpacket),   //          .endofpacket
		.sink5_ready         (crosser_007_out_ready),                 //     sink5.ready
		.sink5_valid         (crosser_007_out_valid),                 //          .valid
		.sink5_channel       (crosser_007_out_channel),               //          .channel
		.sink5_data          (crosser_007_out_data),                  //          .data
		.sink5_startofpacket (crosser_007_out_startofpacket),         //          .startofpacket
		.sink5_endofpacket   (crosser_007_out_endofpacket),           //          .endofpacket
		.sink6_ready         (crosser_009_out_ready),                 //     sink6.ready
		.sink6_valid         (crosser_009_out_valid),                 //          .valid
		.sink6_channel       (crosser_009_out_channel),               //          .channel
		.sink6_data          (crosser_009_out_data),                  //          .data
		.sink6_startofpacket (crosser_009_out_startofpacket),         //          .startofpacket
		.sink6_endofpacket   (crosser_009_out_endofpacket),           //          .endofpacket
		.sink7_ready         (crosser_011_out_ready),                 //     sink7.ready
		.sink7_valid         (crosser_011_out_valid),                 //          .valid
		.sink7_channel       (crosser_011_out_channel),               //          .channel
		.sink7_data          (crosser_011_out_data),                  //          .data
		.sink7_startofpacket (crosser_011_out_startofpacket),         //          .startofpacket
		.sink7_endofpacket   (crosser_011_out_endofpacket)            //          .endofpacket
	);

	soc_system_cmd_xbar_demux_003 cmd_xbar_demux_003 (
		.clk                (pll_sdram_outclk1_clk),                 //       clk.clk
		.reset              (rst_controller_005_reset_out_reset),    // clk_reset.reset
		.sink_ready         (addr_router_003_src_ready),             //      sink.ready
		.sink_channel       (addr_router_003_src_channel),           //          .channel
		.sink_data          (addr_router_003_src_data),              //          .data
		.sink_startofpacket (addr_router_003_src_startofpacket),     //          .startofpacket
		.sink_endofpacket   (addr_router_003_src_endofpacket),       //          .endofpacket
		.sink_valid         (addr_router_003_src_valid),             //          .valid
		.src0_ready         (cmd_xbar_demux_003_src0_ready),         //      src0.ready
		.src0_valid         (cmd_xbar_demux_003_src0_valid),         //          .valid
		.src0_data          (cmd_xbar_demux_003_src0_data),          //          .data
		.src0_channel       (cmd_xbar_demux_003_src0_channel),       //          .channel
		.src0_startofpacket (cmd_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_003_src0_endofpacket)    //          .endofpacket
	);

	soc_system_cmd_xbar_demux_003 cmd_xbar_demux_004 (
		.clk                (pll_sdram_outclk1_clk),                 //       clk.clk
		.reset              (rst_controller_005_reset_out_reset),    // clk_reset.reset
		.sink_ready         (addr_router_004_src_ready),             //      sink.ready
		.sink_channel       (addr_router_004_src_channel),           //          .channel
		.sink_data          (addr_router_004_src_data),              //          .data
		.sink_startofpacket (addr_router_004_src_startofpacket),     //          .startofpacket
		.sink_endofpacket   (addr_router_004_src_endofpacket),       //          .endofpacket
		.sink_valid         (addr_router_004_src_valid),             //          .valid
		.src0_ready         (cmd_xbar_demux_004_src0_ready),         //      src0.ready
		.src0_valid         (cmd_xbar_demux_004_src0_valid),         //          .valid
		.src0_data          (cmd_xbar_demux_004_src0_data),          //          .data
		.src0_channel       (cmd_xbar_demux_004_src0_channel),       //          .channel
		.src0_startofpacket (cmd_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_004_src0_endofpacket)    //          .endofpacket
	);

	soc_system_cmd_xbar_demux_003 cmd_xbar_demux_005 (
		.clk                (pll_sdram_outclk1_clk),                      //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),         // clk_reset.reset
		.sink_ready         (width_adapter_002_cmd_source_ready),         //      sink.ready
		.sink_channel       (width_adapter_002_cmd_source_channel),       //          .channel
		.sink_data          (width_adapter_002_cmd_source_data),          //          .data
		.sink_startofpacket (width_adapter_002_cmd_source_startofpacket), //          .startofpacket
		.sink_endofpacket   (width_adapter_002_cmd_source_endofpacket),   //          .endofpacket
		.sink_valid         (width_adapter_002_cmd_source_valid),         //          .valid
		.src0_ready         (cmd_xbar_demux_005_src0_ready),              //      src0.ready
		.src0_valid         (cmd_xbar_demux_005_src0_valid),              //          .valid
		.src0_data          (cmd_xbar_demux_005_src0_data),               //          .data
		.src0_channel       (cmd_xbar_demux_005_src0_channel),            //          .channel
		.src0_startofpacket (cmd_xbar_demux_005_src0_startofpacket),      //          .startofpacket
		.src0_endofpacket   (cmd_xbar_demux_005_src0_endofpacket)         //          .endofpacket
	);

	soc_system_cmd_xbar_mux_010 cmd_xbar_mux_010 (
		.clk                 (pll_sdram_outclk1_clk),                 //       clk.clk
		.reset               (rst_controller_001_reset_out_reset),    // clk_reset.reset
		.src_ready           (cmd_xbar_mux_010_src_ready),            //       src.ready
		.src_valid           (cmd_xbar_mux_010_src_valid),            //          .valid
		.src_data            (cmd_xbar_mux_010_src_data),             //          .data
		.src_channel         (cmd_xbar_mux_010_src_channel),          //          .channel
		.src_startofpacket   (cmd_xbar_mux_010_src_startofpacket),    //          .startofpacket
		.src_endofpacket     (cmd_xbar_mux_010_src_endofpacket),      //          .endofpacket
		.sink0_ready         (cmd_xbar_demux_003_src0_ready),         //     sink0.ready
		.sink0_valid         (cmd_xbar_demux_003_src0_valid),         //          .valid
		.sink0_channel       (cmd_xbar_demux_003_src0_channel),       //          .channel
		.sink0_data          (cmd_xbar_demux_003_src0_data),          //          .data
		.sink0_startofpacket (cmd_xbar_demux_003_src0_startofpacket), //          .startofpacket
		.sink0_endofpacket   (cmd_xbar_demux_003_src0_endofpacket),   //          .endofpacket
		.sink1_ready         (cmd_xbar_demux_004_src0_ready),         //     sink1.ready
		.sink1_valid         (cmd_xbar_demux_004_src0_valid),         //          .valid
		.sink1_channel       (cmd_xbar_demux_004_src0_channel),       //          .channel
		.sink1_data          (cmd_xbar_demux_004_src0_data),          //          .data
		.sink1_startofpacket (cmd_xbar_demux_004_src0_startofpacket), //          .startofpacket
		.sink1_endofpacket   (cmd_xbar_demux_004_src0_endofpacket),   //          .endofpacket
		.sink2_ready         (cmd_xbar_demux_005_src0_ready),         //     sink2.ready
		.sink2_valid         (cmd_xbar_demux_005_src0_valid),         //          .valid
		.sink2_channel       (cmd_xbar_demux_005_src0_channel),       //          .channel
		.sink2_data          (cmd_xbar_demux_005_src0_data),          //          .data
		.sink2_startofpacket (cmd_xbar_demux_005_src0_startofpacket), //          .startofpacket
		.sink2_endofpacket   (cmd_xbar_demux_005_src0_endofpacket)    //          .endofpacket
	);

	soc_system_rsp_xbar_demux_010 rsp_xbar_demux_010 (
		.clk                (pll_sdram_outclk1_clk),                      //       clk.clk
		.reset              (rst_controller_001_reset_out_reset),         // clk_reset.reset
		.sink_ready         (width_adapter_003_rsp_source_ready),         //      sink.ready
		.sink_channel       (width_adapter_003_rsp_source_channel),       //          .channel
		.sink_data          (width_adapter_003_rsp_source_data),          //          .data
		.sink_startofpacket (width_adapter_003_rsp_source_startofpacket), //          .startofpacket
		.sink_endofpacket   (width_adapter_003_rsp_source_endofpacket),   //          .endofpacket
		.sink_valid         (width_adapter_003_rsp_source_valid),         //          .valid
		.src0_ready         (rsp_xbar_demux_010_src0_ready),              //      src0.ready
		.src0_valid         (rsp_xbar_demux_010_src0_valid),              //          .valid
		.src0_data          (rsp_xbar_demux_010_src0_data),               //          .data
		.src0_channel       (rsp_xbar_demux_010_src0_channel),            //          .channel
		.src0_startofpacket (rsp_xbar_demux_010_src0_startofpacket),      //          .startofpacket
		.src0_endofpacket   (rsp_xbar_demux_010_src0_endofpacket),        //          .endofpacket
		.src1_ready         (rsp_xbar_demux_010_src1_ready),              //      src1.ready
		.src1_valid         (rsp_xbar_demux_010_src1_valid),              //          .valid
		.src1_data          (rsp_xbar_demux_010_src1_data),               //          .data
		.src1_channel       (rsp_xbar_demux_010_src1_channel),            //          .channel
		.src1_startofpacket (rsp_xbar_demux_010_src1_startofpacket),      //          .startofpacket
		.src1_endofpacket   (rsp_xbar_demux_010_src1_endofpacket),        //          .endofpacket
		.src2_ready         (rsp_xbar_demux_010_src2_ready),              //      src2.ready
		.src2_valid         (rsp_xbar_demux_010_src2_valid),              //          .valid
		.src2_data          (rsp_xbar_demux_010_src2_data),               //          .data
		.src2_channel       (rsp_xbar_demux_010_src2_channel),            //          .channel
		.src2_startofpacket (rsp_xbar_demux_010_src2_startofpacket),      //          .startofpacket
		.src2_endofpacket   (rsp_xbar_demux_010_src2_endofpacket)         //          .endofpacket
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (113),
		.BITS_PER_SYMBOL     (113),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (8),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser (
		.in_clk            (clk_clk),                               //        in_clk.clk
		.in_reset          (rst_controller_004_reset_out_reset),    //  in_clk_reset.reset
		.out_clk           (pll_stream_outclk1_clk),                //       out_clk.clk
		.out_reset         (rst_controller_002_reset_out_reset),    // out_clk_reset.reset
		.in_ready          (cmd_xbar_demux_001_src5_ready),         //            in.ready
		.in_valid          (cmd_xbar_demux_001_src5_valid),         //              .valid
		.in_startofpacket  (cmd_xbar_demux_001_src5_startofpacket), //              .startofpacket
		.in_endofpacket    (cmd_xbar_demux_001_src5_endofpacket),   //              .endofpacket
		.in_channel        (cmd_xbar_demux_001_src5_channel),       //              .channel
		.in_data           (cmd_xbar_demux_001_src5_data),          //              .data
		.out_ready         (crosser_out_ready),                     //           out.ready
		.out_valid         (crosser_out_valid),                     //              .valid
		.out_startofpacket (crosser_out_startofpacket),             //              .startofpacket
		.out_endofpacket   (crosser_out_endofpacket),               //              .endofpacket
		.out_channel       (crosser_out_channel),                   //              .channel
		.out_data          (crosser_out_data),                      //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (113),
		.BITS_PER_SYMBOL     (113),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (8),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_001 (
		.in_clk            (clk_clk),                               //        in_clk.clk
		.in_reset          (rst_controller_004_reset_out_reset),    //  in_clk_reset.reset
		.out_clk           (pll_stream_outclk1_clk),                //       out_clk.clk
		.out_reset         (rst_controller_002_reset_out_reset),    // out_clk_reset.reset
		.in_ready          (cmd_xbar_demux_001_src6_ready),         //            in.ready
		.in_valid          (cmd_xbar_demux_001_src6_valid),         //              .valid
		.in_startofpacket  (cmd_xbar_demux_001_src6_startofpacket), //              .startofpacket
		.in_endofpacket    (cmd_xbar_demux_001_src6_endofpacket),   //              .endofpacket
		.in_channel        (cmd_xbar_demux_001_src6_channel),       //              .channel
		.in_data           (cmd_xbar_demux_001_src6_data),          //              .data
		.out_ready         (crosser_001_out_ready),                 //           out.ready
		.out_valid         (crosser_001_out_valid),                 //              .valid
		.out_startofpacket (crosser_001_out_startofpacket),         //              .startofpacket
		.out_endofpacket   (crosser_001_out_endofpacket),           //              .endofpacket
		.out_channel       (crosser_001_out_channel),               //              .channel
		.out_data          (crosser_001_out_data),                  //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (113),
		.BITS_PER_SYMBOL     (113),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (8),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_002 (
		.in_clk            (clk_clk),                               //        in_clk.clk
		.in_reset          (rst_controller_004_reset_out_reset),    //  in_clk_reset.reset
		.out_clk           (pll_audio_outclk0_clk),                 //       out_clk.clk
		.out_reset         (rst_controller_003_reset_out_reset),    // out_clk_reset.reset
		.in_ready          (cmd_xbar_demux_001_src7_ready),         //            in.ready
		.in_valid          (cmd_xbar_demux_001_src7_valid),         //              .valid
		.in_startofpacket  (cmd_xbar_demux_001_src7_startofpacket), //              .startofpacket
		.in_endofpacket    (cmd_xbar_demux_001_src7_endofpacket),   //              .endofpacket
		.in_channel        (cmd_xbar_demux_001_src7_channel),       //              .channel
		.in_data           (cmd_xbar_demux_001_src7_data),          //              .data
		.out_ready         (crosser_002_out_ready),                 //           out.ready
		.out_valid         (crosser_002_out_valid),                 //              .valid
		.out_startofpacket (crosser_002_out_startofpacket),         //              .startofpacket
		.out_endofpacket   (crosser_002_out_endofpacket),           //              .endofpacket
		.out_channel       (crosser_002_out_channel),               //              .channel
		.out_data          (crosser_002_out_data),                  //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (113),
		.BITS_PER_SYMBOL     (113),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (8),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_003 (
		.in_clk            (clk_clk),                               //        in_clk.clk
		.in_reset          (rst_controller_004_reset_out_reset),    //  in_clk_reset.reset
		.out_clk           (pll_stream_outclk1_clk),                //       out_clk.clk
		.out_reset         (rst_controller_002_reset_out_reset),    // out_clk_reset.reset
		.in_ready          (cmd_xbar_demux_002_src5_ready),         //            in.ready
		.in_valid          (cmd_xbar_demux_002_src5_valid),         //              .valid
		.in_startofpacket  (cmd_xbar_demux_002_src5_startofpacket), //              .startofpacket
		.in_endofpacket    (cmd_xbar_demux_002_src5_endofpacket),   //              .endofpacket
		.in_channel        (cmd_xbar_demux_002_src5_channel),       //              .channel
		.in_data           (cmd_xbar_demux_002_src5_data),          //              .data
		.out_ready         (crosser_003_out_ready),                 //           out.ready
		.out_valid         (crosser_003_out_valid),                 //              .valid
		.out_startofpacket (crosser_003_out_startofpacket),         //              .startofpacket
		.out_endofpacket   (crosser_003_out_endofpacket),           //              .endofpacket
		.out_channel       (crosser_003_out_channel),               //              .channel
		.out_data          (crosser_003_out_data),                  //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (113),
		.BITS_PER_SYMBOL     (113),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (8),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_004 (
		.in_clk            (clk_clk),                               //        in_clk.clk
		.in_reset          (rst_controller_004_reset_out_reset),    //  in_clk_reset.reset
		.out_clk           (pll_stream_outclk1_clk),                //       out_clk.clk
		.out_reset         (rst_controller_002_reset_out_reset),    // out_clk_reset.reset
		.in_ready          (cmd_xbar_demux_002_src6_ready),         //            in.ready
		.in_valid          (cmd_xbar_demux_002_src6_valid),         //              .valid
		.in_startofpacket  (cmd_xbar_demux_002_src6_startofpacket), //              .startofpacket
		.in_endofpacket    (cmd_xbar_demux_002_src6_endofpacket),   //              .endofpacket
		.in_channel        (cmd_xbar_demux_002_src6_channel),       //              .channel
		.in_data           (cmd_xbar_demux_002_src6_data),          //              .data
		.out_ready         (crosser_004_out_ready),                 //           out.ready
		.out_valid         (crosser_004_out_valid),                 //              .valid
		.out_startofpacket (crosser_004_out_startofpacket),         //              .startofpacket
		.out_endofpacket   (crosser_004_out_endofpacket),           //              .endofpacket
		.out_channel       (crosser_004_out_channel),               //              .channel
		.out_data          (crosser_004_out_data),                  //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (113),
		.BITS_PER_SYMBOL     (113),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (8),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_005 (
		.in_clk            (clk_clk),                               //        in_clk.clk
		.in_reset          (rst_controller_004_reset_out_reset),    //  in_clk_reset.reset
		.out_clk           (pll_audio_outclk0_clk),                 //       out_clk.clk
		.out_reset         (rst_controller_003_reset_out_reset),    // out_clk_reset.reset
		.in_ready          (cmd_xbar_demux_002_src7_ready),         //            in.ready
		.in_valid          (cmd_xbar_demux_002_src7_valid),         //              .valid
		.in_startofpacket  (cmd_xbar_demux_002_src7_startofpacket), //              .startofpacket
		.in_endofpacket    (cmd_xbar_demux_002_src7_endofpacket),   //              .endofpacket
		.in_channel        (cmd_xbar_demux_002_src7_channel),       //              .channel
		.in_data           (cmd_xbar_demux_002_src7_data),          //              .data
		.out_ready         (crosser_005_out_ready),                 //           out.ready
		.out_valid         (crosser_005_out_valid),                 //              .valid
		.out_startofpacket (crosser_005_out_startofpacket),         //              .startofpacket
		.out_endofpacket   (crosser_005_out_endofpacket),           //              .endofpacket
		.out_channel       (crosser_005_out_channel),               //              .channel
		.out_data          (crosser_005_out_data),                  //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (113),
		.BITS_PER_SYMBOL     (113),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (8),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_006 (
		.in_clk            (pll_stream_outclk1_clk),                //        in_clk.clk
		.in_reset          (rst_controller_002_reset_out_reset),    //  in_clk_reset.reset
		.out_clk           (clk_clk),                               //       out_clk.clk
		.out_reset         (rst_controller_004_reset_out_reset),    // out_clk_reset.reset
		.in_ready          (rsp_xbar_demux_007_src0_ready),         //            in.ready
		.in_valid          (rsp_xbar_demux_007_src0_valid),         //              .valid
		.in_startofpacket  (rsp_xbar_demux_007_src0_startofpacket), //              .startofpacket
		.in_endofpacket    (rsp_xbar_demux_007_src0_endofpacket),   //              .endofpacket
		.in_channel        (rsp_xbar_demux_007_src0_channel),       //              .channel
		.in_data           (rsp_xbar_demux_007_src0_data),          //              .data
		.out_ready         (crosser_006_out_ready),                 //           out.ready
		.out_valid         (crosser_006_out_valid),                 //              .valid
		.out_startofpacket (crosser_006_out_startofpacket),         //              .startofpacket
		.out_endofpacket   (crosser_006_out_endofpacket),           //              .endofpacket
		.out_channel       (crosser_006_out_channel),               //              .channel
		.out_data          (crosser_006_out_data),                  //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (113),
		.BITS_PER_SYMBOL     (113),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (8),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_007 (
		.in_clk            (pll_stream_outclk1_clk),                //        in_clk.clk
		.in_reset          (rst_controller_002_reset_out_reset),    //  in_clk_reset.reset
		.out_clk           (clk_clk),                               //       out_clk.clk
		.out_reset         (rst_controller_004_reset_out_reset),    // out_clk_reset.reset
		.in_ready          (rsp_xbar_demux_007_src1_ready),         //            in.ready
		.in_valid          (rsp_xbar_demux_007_src1_valid),         //              .valid
		.in_startofpacket  (rsp_xbar_demux_007_src1_startofpacket), //              .startofpacket
		.in_endofpacket    (rsp_xbar_demux_007_src1_endofpacket),   //              .endofpacket
		.in_channel        (rsp_xbar_demux_007_src1_channel),       //              .channel
		.in_data           (rsp_xbar_demux_007_src1_data),          //              .data
		.out_ready         (crosser_007_out_ready),                 //           out.ready
		.out_valid         (crosser_007_out_valid),                 //              .valid
		.out_startofpacket (crosser_007_out_startofpacket),         //              .startofpacket
		.out_endofpacket   (crosser_007_out_endofpacket),           //              .endofpacket
		.out_channel       (crosser_007_out_channel),               //              .channel
		.out_data          (crosser_007_out_data),                  //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (113),
		.BITS_PER_SYMBOL     (113),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (8),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_008 (
		.in_clk            (pll_stream_outclk1_clk),                //        in_clk.clk
		.in_reset          (rst_controller_002_reset_out_reset),    //  in_clk_reset.reset
		.out_clk           (clk_clk),                               //       out_clk.clk
		.out_reset         (rst_controller_004_reset_out_reset),    // out_clk_reset.reset
		.in_ready          (rsp_xbar_demux_008_src0_ready),         //            in.ready
		.in_valid          (rsp_xbar_demux_008_src0_valid),         //              .valid
		.in_startofpacket  (rsp_xbar_demux_008_src0_startofpacket), //              .startofpacket
		.in_endofpacket    (rsp_xbar_demux_008_src0_endofpacket),   //              .endofpacket
		.in_channel        (rsp_xbar_demux_008_src0_channel),       //              .channel
		.in_data           (rsp_xbar_demux_008_src0_data),          //              .data
		.out_ready         (crosser_008_out_ready),                 //           out.ready
		.out_valid         (crosser_008_out_valid),                 //              .valid
		.out_startofpacket (crosser_008_out_startofpacket),         //              .startofpacket
		.out_endofpacket   (crosser_008_out_endofpacket),           //              .endofpacket
		.out_channel       (crosser_008_out_channel),               //              .channel
		.out_data          (crosser_008_out_data),                  //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (113),
		.BITS_PER_SYMBOL     (113),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (8),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_009 (
		.in_clk            (pll_stream_outclk1_clk),                //        in_clk.clk
		.in_reset          (rst_controller_002_reset_out_reset),    //  in_clk_reset.reset
		.out_clk           (clk_clk),                               //       out_clk.clk
		.out_reset         (rst_controller_004_reset_out_reset),    // out_clk_reset.reset
		.in_ready          (rsp_xbar_demux_008_src1_ready),         //            in.ready
		.in_valid          (rsp_xbar_demux_008_src1_valid),         //              .valid
		.in_startofpacket  (rsp_xbar_demux_008_src1_startofpacket), //              .startofpacket
		.in_endofpacket    (rsp_xbar_demux_008_src1_endofpacket),   //              .endofpacket
		.in_channel        (rsp_xbar_demux_008_src1_channel),       //              .channel
		.in_data           (rsp_xbar_demux_008_src1_data),          //              .data
		.out_ready         (crosser_009_out_ready),                 //           out.ready
		.out_valid         (crosser_009_out_valid),                 //              .valid
		.out_startofpacket (crosser_009_out_startofpacket),         //              .startofpacket
		.out_endofpacket   (crosser_009_out_endofpacket),           //              .endofpacket
		.out_channel       (crosser_009_out_channel),               //              .channel
		.out_data          (crosser_009_out_data),                  //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (113),
		.BITS_PER_SYMBOL     (113),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (8),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_010 (
		.in_clk            (pll_audio_outclk0_clk),                 //        in_clk.clk
		.in_reset          (rst_controller_003_reset_out_reset),    //  in_clk_reset.reset
		.out_clk           (clk_clk),                               //       out_clk.clk
		.out_reset         (rst_controller_004_reset_out_reset),    // out_clk_reset.reset
		.in_ready          (rsp_xbar_demux_009_src0_ready),         //            in.ready
		.in_valid          (rsp_xbar_demux_009_src0_valid),         //              .valid
		.in_startofpacket  (rsp_xbar_demux_009_src0_startofpacket), //              .startofpacket
		.in_endofpacket    (rsp_xbar_demux_009_src0_endofpacket),   //              .endofpacket
		.in_channel        (rsp_xbar_demux_009_src0_channel),       //              .channel
		.in_data           (rsp_xbar_demux_009_src0_data),          //              .data
		.out_ready         (crosser_010_out_ready),                 //           out.ready
		.out_valid         (crosser_010_out_valid),                 //              .valid
		.out_startofpacket (crosser_010_out_startofpacket),         //              .startofpacket
		.out_endofpacket   (crosser_010_out_endofpacket),           //              .endofpacket
		.out_channel       (crosser_010_out_channel),               //              .channel
		.out_data          (crosser_010_out_data),                  //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	altera_avalon_st_handshake_clock_crosser #(
		.DATA_WIDTH          (113),
		.BITS_PER_SYMBOL     (113),
		.USE_PACKETS         (1),
		.USE_CHANNEL         (1),
		.CHANNEL_WIDTH       (8),
		.USE_ERROR           (0),
		.ERROR_WIDTH         (1),
		.VALID_SYNC_DEPTH    (2),
		.READY_SYNC_DEPTH    (2),
		.USE_OUTPUT_PIPELINE (0)
	) crosser_011 (
		.in_clk            (pll_audio_outclk0_clk),                 //        in_clk.clk
		.in_reset          (rst_controller_003_reset_out_reset),    //  in_clk_reset.reset
		.out_clk           (clk_clk),                               //       out_clk.clk
		.out_reset         (rst_controller_004_reset_out_reset),    // out_clk_reset.reset
		.in_ready          (rsp_xbar_demux_009_src1_ready),         //            in.ready
		.in_valid          (rsp_xbar_demux_009_src1_valid),         //              .valid
		.in_startofpacket  (rsp_xbar_demux_009_src1_startofpacket), //              .startofpacket
		.in_endofpacket    (rsp_xbar_demux_009_src1_endofpacket),   //              .endofpacket
		.in_channel        (rsp_xbar_demux_009_src1_channel),       //              .channel
		.in_data           (rsp_xbar_demux_009_src1_data),          //              .data
		.out_ready         (crosser_011_out_ready),                 //           out.ready
		.out_valid         (crosser_011_out_valid),                 //              .valid
		.out_startofpacket (crosser_011_out_startofpacket),         //              .startofpacket
		.out_endofpacket   (crosser_011_out_endofpacket),           //              .endofpacket
		.out_channel       (crosser_011_out_channel),               //              .channel
		.out_data          (crosser_011_out_data),                  //              .data
		.in_empty          (1'b0),                                  //   (terminated)
		.in_error          (1'b0),                                  //   (terminated)
		.out_empty         (),                                      //   (terminated)
		.out_error         ()                                       //   (terminated)
	);

	soc_system_irq_mapper irq_mapper (
		.clk           (),                         //       clk.clk
		.reset         (),                         // clk_reset.reset
		.receiver0_irq (irq_mapper_receiver0_irq), // receiver0.irq
		.receiver1_irq (irq_mapper_receiver1_irq), // receiver1.irq
		.receiver2_irq (irq_mapper_receiver2_irq), // receiver2.irq
		.sender_irq    (hps_0_f2h_irq0_irq)        //    sender.irq
	);

	soc_system_irq_mapper_001 irq_mapper_001 (
		.clk        (),                   //       clk.clk
		.reset      (),                   // clk_reset.reset
		.sender_irq (hps_0_f2h_irq1_irq)  //    sender.irq
	);

	soc_system_avalon_st_adapter #(
		.inBitsPerSymbol (8),
		.inUsePackets    (1),
		.inDataWidth     (24),
		.inChannelWidth  (0),
		.inErrorWidth    (0),
		.inUseEmptyPort  (1),
		.inUseValid      (1),
		.inUseReady      (1),
		.inReadyLatency  (1),
		.outDataWidth    (24),
		.outChannelWidth (0),
		.outErrorWidth   (0),
		.outUseEmptyPort (0),
		.outUseValid     (1),
		.outUseReady     (1),
		.outReadyLatency (0)
	) avalon_st_adapter (
		.in_clk_0_clk        (pll_stream_outclk1_clk),                // in_clk_0.clk
		.in_rst_0_reset      (rst_controller_002_reset_out_reset),    // in_rst_0.reset
		.in_0_ready          (log_generate_0_dout_ready),             //     in_0.ready
		.in_0_valid          (log_generate_0_dout_valid),             //         .valid
		.in_0_data           (log_generate_0_dout_data),              //         .data
		.in_0_startofpacket  (log_generate_0_dout_startofpacket),     //         .startofpacket
		.in_0_endofpacket    (log_generate_0_dout_endofpacket),       //         .endofpacket
		.in_0_empty          (log_generate_0_dout_empty),             //         .empty
		.out_0_ready         (avalon_st_adapter_out_0_ready),         //    out_0.ready
		.out_0_valid         (avalon_st_adapter_out_0_valid),         //         .valid
		.out_0_data          (avalon_st_adapter_out_0_data),          //         .data
		.out_0_startofpacket (avalon_st_adapter_out_0_startofpacket), //         .startofpacket
		.out_0_endofpacket   (avalon_st_adapter_out_0_endofpacket)    //         .endofpacket
	);

endmodule
