��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%�����d^S$�0���<SG���0}�q�hS���.o�o�X{R�?9�x��ּ�@�����Y�v.'1t��>�1M=�\,�i�R5V[d�
�����@Xk���Fq���$Z�u�չ���J 	��Ǐ�J;a��^��?�o{̛����
�Fb�G�f��ۤ`U���oȚ�ufJ���g>U�;0�)�[��[\C٧��Wi���a͟��aoOL���D���Kj�h�4?��n%NE:Yi����Ǟ�H� �a�C�����c�&�|�ۣ"�6����=a�BT7�](���~�՜�l�ܞ&�f:XΕ�B�:�,=��Q9{Våi��}Q(:&o`�G�5�e^�5���3�n���� �c��1!Hz�'�<~23�@��[��"�{�U~�*+6��Pn����N:�|���p�\.W5�?����	r�{��9c�g��;����������>�ߴ0$Ǿ��Պ~�Q<X��Ԙ[A/ԗ���lZ��Q���ݾ�60:p�+���2��|��a��������~wα�=|s����g�c!�X�o��m���RPI�-��Q��gL��.�� ��wv *���	q�c,*�`
��<�r)�m� ��v������Ӝ8��B9+��c,U]���L٢zvK�C$��\�J]��K�]t��z�hAˡͶ� <�kM���8�Y�nX;�u�AM���݇*y)�I�=�݂ᯢI��a���A�)#j��(��_�|��	2S��G[�s�J�L���m��ݼ�mH�̓��Z�O���%F�Y��c���I�cAIʸ�(^�ʷ��}Im~P�	��MP�Y��'�ϧJj���<&8�][�
T<�����`_É���g�Y�`����YjML��J������%L�����n?��)�`.��7�B8�˯�{e{�M .��|s�<�%�`ф���8P"�dm��Cpl5���pK��+᠙�F��#+ֆW�
�>*ɻ�Y�����bc���f��sX-�����zn��������өC�m`��+)]v���=�
���f�a4{�y��'K,r�8e����s�)��b�,����U�8��n�P�ˊGt�"b~ڐ�.�D<��Z;�������7��y�z�0�eA�`&�q9��R�	�5���|��WB���b�ݢ�a�g�K���h� ����\���o�p<�//O�P��x��BN�64n�P��[7��Å�pBY��
1*VU��>o�q2�M����ʷ�iT�U���i�3.⠷���g��L��9�n�����J���;��y���4o;���^������G�����"&�A�����S�D����i.DV��N��hF7�^�ף�"],��Q���6Dv�Ֆ�߮z��~R��?���MaF��'g����tĴ����2 �	�e�U�*L���'x�������f/�����^\�&�dP�w_�:k�L��^6-�z��IpnT#��E�jF�n`���	�P*O����XMeX<14	'�d>��LϽo}��scƾ4��Cpd�Җ�r�;xdA��70B_Ku(O�y�z�Dn���C��~�����R�m� ��Z���>>�V��Qb���p��_��J>��'�$rZ����.��>�R��R�
�e\h��-!U��r8�&Hk���߁����p1��|���0�jٴ݇N=�#(�� J�Y�ӿE��he_����4��b�
�''̨� �?�gA����>	Z��ҶW��,�c��4���V�j��<(�-�	m9IC�<��j*�x�K���\;XKXS��X�/I��Z[x���A��񟯺S�T9	b2�� �B����w�lE�*y��x�)���ɞS�.�I���YNl��!T��v��v|��"���kT���f+��)��`�$I|�^�5G1&x������)�^� v���ً�xo�{Tw �l���p#�+����)�
���͗�N��'wmNμ�X�'S�2;��J�r� �����Q�Qj_��d^kmd�9�H����&�|���LE�t��%�]k-���t�e[�>�=aP�r��E��-
�r���$����^�ZЁlx��]��遵e$����ʈ66m����x��<��ޫ�R>���6���h����^�űW�%�
s�_#w�5��<�i��	\��?��O��ωF�{�"�M�ڬ����`�OC0��"\�u��F�I64D1�S�-Wm�KT��YloR��8ȴ>�z2�b�o]�g(;u�2V�^�~xd���&3��8(N����|�v�Ѝ9���:3�bܺ%�y�	$��/�r�䴇��㣋(
�/96ݲ��)�!���߈@��"e�0B�w�3-�@��e�N*���d�}`��ND�����H�����(��M�@�<f��e��P��$��p��L����yJ�]\�������I_�fO~bU�}'�Ψ%�Ֆ9;�(yV��1T����Ni������J�1���"�n��v�vԺbU��W��+����
9]����Ψq�E�޵��(V?��d���J4x	T;D���v��O�;J@��\�x�o��Vǂ��X�����P��h.�����/�<sI�����ngM��N��>�����Ы����RZ�㞸�l#~��ܓR=ZXj�VO,/��H���>�2M��+�Ф�Ma����C6+������,���,r�&��֎���:�sg��,���fP����ڪv��)�T�@�h��V,O��!�_Eg�'�������R͉�'^%��?Z"���$��̈́�2�������_nj����ţ>��9&�\�K��
{���m��s��HI�F�
*�����B_a����� ��PG����E~ǋ��+�Z�\s� �ܺx�� Y���J�/���D÷��*���k����g�JL�3�4�.$"M����3���{|pt%�x�-��1x�y��tn�GP�j�dV��p~n�I�'h�`j�,M������؀(\�{+[Z�e
R�tj,˿����]'�vD�ky�9}�w@��1�(*D�@�����w����+[�e~/�Q0���>&g!s��"w�L'�S�C�w����\�W
�/Y�Ƌ�'܄'�9�$��;�'�e"�GW	�ng2�O[�p���,� XCt�˾t.�|.��g ���'�����
Crk�FS9�dx�®o�<	��d�-,T�:�&N�*YB�C����&]���Z�mmLw���iѠ�ux�T��X�?�2�L��E4���ѻո�pHK���>�u�gۿh�Вx�W}�^����a<���·O+�42��g�x3yg���4��J�������X&g�-����fa�G�v��.kV2�A)�32�`�O����Ϡ��a������6�_�QM;���pXP�e�� Gn?Q��2����d��Y��[��A��N<� �� ��I�d��cvW��v�bE�����y.;��"�Ԓ�2 �.��E1jGz���`�3�m���f�����<k����oǧ��b���w�\�� ݿy�����(Jb8���Bo�f�:�R�5������dG��d:*@���ܹ��qB�'>l��qT<����X�#S��h��P�'籹�/s�;�!"�3ӿJ�%	V�f��Q�2]����?eNO���k<o� 6p|�6���?����J��]_I�R���<�U���5�\�z�L�A_����(�DZm�p~��c��(�K���E�?&�}���k�il�����g�:5ԍ<D��K84�F�D���N{��P7����].�/h%;|�+h���ܨ"�ZC65pC��,��4����cK��q��i�E�'&yȻ�%?kC��ݶ�6A�1̀]�ע�V��
���%��_�N�|�Z����SE�����gA�1o�0rk���dm�K7�2����F�X������7�6���y"{��]��7��R�
9룝#��w�"v;����� Gw�&}�àa&Z���0�ؑ/�E;q'"�Z�Ǖe2��v��uuS��91W/��[.ʵK�Nj,��V�5ƴ\8��,2Td�g�9Ӈ��V���Mj�̇ؿ�Z	�&*zj0��NEל>qS�� ��؟����#e�w$���좚2J\P������~�Y����a��A����#t��w�Ⱥ�9������Xk#\�eJѸ���@����߃{��t�d'?��o�<Z�;�?��o|\N��>8'��S鷵=�TD�����2���9��N�ӰH�����&��9p%�(������ y�~�2U���[�q���1��k�T�y����ڡ���ʳ Q��K~Eov &1��F��ϴ��R|j��v�F�r�
�`�k�zf��� ���D�D+��	�&�(�h�1lV_�µ��H�,����!�ꚽD�Iˀ7/���F���8��,G��E����7ԝ2��|ˁ�e�k�����@�r�E_�ҝ�k��y����n���{&� !�`aEp�H��3�޸I�Or�^�v'�r�B����I6)�a��F �,W���*�� �z�Dd�go�|�L-s�q��{�v�gˌ�q5�Ka� �y섳9�Zr+&�.Z�rj�'�a��&:��à����
�O��вjI�G[=)QVM�H�l20�Rr$�4�	O2���D��"���'̭�X�
u������\�l����QeA'R�	h��Q�ػ'�=���p��S�"�5��DM�����&��-o3�@<�j����:O��1���{�3�ZЪf�]g�������������I�m���(�I�z
&�9r�!XJ�h&�@|�>�l8�����f���#�V��%�]���A��y�Z��U�WAB�&
IS�\��0I,ʥ��f���yW��e�PiUY�-�GL'L]\�yΈ�1s�e ���~(��#�Z��B�m^����3cP��}��I�ٌ�XDY+!�������Y����#��Q���u�}B��/R������sKAx=kW�G�Yfu�ط��8��c�{�ڗ�y�-V�8>�����6��Z���h���2ִ�X�&^�.oM��&��?4�q�rc��N��^�4��Q�KZI����(#&ya=����,o�3�m�������F�mf�,��J��k��5�����N�^�J#��s��Dh��2�Nl��Ž��s��3�.����b:�˛�L̖�.��*<��V�}�j����C�$��5(D�>$�xj]���V䅞�)�yv�%�mhZ,V���t	ަ�0��h��tY�d�&�oE�.�.�����
��j���:-?m`����!���'wHD8ОR,�~�j/��] ���@�'4��PX�˦�3J����o�:Rpb^��K�����	���Ea"�����w��ܗ���Ke5
�͢��-�����L��z(ͣ��kM�z���ZV�s�C���%��~6q�d#����\N���+��O�z>���'s*�o�9 ^Nc���D´+,���� �&�2� �x�ZL�DNJ�rkS�8�P���e�ra*	��+z�o=u�8#9���;<_!�۟S�S���ʣ"��p�� p}����|���!@��s�L����j��:b�j��d��X�QQE�HtG����X�oyI�c��۷��B��j�3��(��d�|w%'�Z��K�w���5E���%N�NG�^���l�r���nWL����m^c�X�y�v����sR>��&���A9I� �R���g��h���-{7I���TL����D���f��[���.1�1����/�+ۏ��A����.���PpK� 	�ٝS-�_ �r�l5N�}Α���'���Mu�u���F�R�"��8ղ�x
���H
?�؆'���Q܊�xZ�<⟖�ؠ�O��rM�zns��r��H>�I�C�}\���Fg6j��\_<J�ƶ�8����Bĵ�B�=Z�v��]��w�wSJ���p揩���6[a�ńa��-���4f8��S�4THd���9UҔf���6[�|g�m�T�`� �o�7��b7��>�� ���:���b�	����K0���Z�w��������l���H�|����4���V4=E�g����I���M��r�_���n{A$������'�h�yr����n��N4���L�z�� ���[���@Q�V'[P{�`od����F��JV܁o���c�JD{�q�a���	�z��M��w@��Ų�yvǨ�j����'��W ��4]����)pƈz����DS�&]�#���u=bb̾������G[\l`CS���j���Y�w���wX�G�U�+/�)� U��l$��f
���*,����9.,�'7��*H�8D��y��F29�v>�+�;����$��>�ЃI�VRG�����x�n�{�SR_0U�� ���ط8.�Z�S s��іV��$�4�%�e�aP��+>���"Q�R'(c��b�z��?�O�t���l`.�0�_�\%���1�s�>��щ_���k��4�0N�x��Ḋ݂��AqSjq�	�Q>R:��A�ܼ�_'�󇟑�*'����s7#��^�����s�CX}�SyL��;?u����$�_�=ڃ���mT[�C��*��Dk�Q]�8ۖ[��e�;�)ĳ:wcvɭ���?WȐY��d�v�Wݶ4�HbĲ y�i����l�ޏL��>[I����j���[#���ڒһ̗�x��&
n:�7�yp������x`���N����_;��� �4)���e�/�bL�aA�ڑ�_~��g|dKu��"���0�B��lXO�ۨX	�yA�߯���[���eH��J�=��R=f�Њ?����iƍ��KE�~t����>�_Ā�{����:��\K�,Y��w�NB��n&�H4�`��"�(�D�Z�*x�" *=1v�H�k�u�ZU):m�a)��輤V"��k���L����F��nb=R��;,��aᙞ�����먼���x��ȍ��~)L�O�H-�ΣkӶgH��q�f��j1�>k�|�-�/�k��O�5c���2�`$����q_��:2�.��C�	s�?�"��A�g
FІN�In�C����a,�1����3aD$��������D+�<�XNx2g���5�/�Ӷ#�է��\�	��'�[���a�O9lCa��Qyi��y�:���|�`���h��OL��HK0K�^�k�G[�slB5�m�-_~��K�s�8��.���خ�;S�2Cbɬ=���]0�paɰȥv�{t�Z�M1j�k��Dlg�=[Iz�,�%L���0!6���m��򔰛)�U�j�� 6uY8�S�q����t"�\�Up��r�g�\�hjT�B����K%���������Ⰻyў�\�I��7Z�&ƶ����ҏ�ђc�i�Dd�6���DY����"��[�h+2M��#pW8���6I�)�(d ��k|TU7%��#�V�LOj
����~�T����Bn���O� yT����$����	�D�W�Ϫ9�3�nC}��9%ATj���kb#nGc�[�괙/w.�fɩnu��͐^��@�v*�y?��6꿠MZf��Id��_I�ŏ�	�`W�2� !�w� \���RlY����ɮ�N��?4��Y���0�~�h%w�-�o���ݖz���XEc	��ip�݇��s��J�l	V?/��l���p�k�Q��C'��vD�� ��wޅ�+Ze'�&���?�j�a���*`F�l[����p_m݁
�n����\�@�yK�5� АV�}����9�#�h 5[Q�l���]H} uO�����\Zϓ�	u�`���"���w�+��lk�ޖ���_�\g�+�r�(W||�>{���Ş��\?xv���r�Zi��ap�v3%�8w�Z��pIbm��^qeI�~��w�-7���ś��K*&����U��ޮf���L������wVǼށ��"��!���a��JE��ހ��x�{C�Ŋ�(����&?�Z*�=�G��͎������A� �5�,�rg�O��G�,��ِ;;Y	���O�c���ɗ��B~�t�M0Ϟ_��O�9� �~�n*^�ҍ��L	�X�F�z?B(�a�SW��w,�&.%����j �����H��l�=�b"�0��ӱ{��}u�l^ba.���]�� ��S�#�\EJx{�������3f�u����Q�����6��U����Y�J�M퀿|_��ѐ�~6�2.⏯KS�Sn���Vv�B���r��'���s�U`#��mb�XL���N�r�T4J'L����n���#c�Do�h�
wG���|[���?i]����x�f"�#K�Đ�d���Vz�,��~!� :5˄*�������Uh�ƪ����<�Z5o��>���_]��~�K���.N ~)���:�H{7��h�[��,�+n���,�(����@X3VajhBO	p�W���dig������*Y�v�a�#tI2�'k�\I�J8J�3��3�����C眢R6L��gZ�-	g�.�~�gT�tb�+K�/�!�9�N-��`���?��7��K�ߌ�Tk�$i�I�%���a�}��;����.Oq��'�d�ov8��˥)!��a���z�p�V�M?Ii�k-*6��`i��������~�e\6�d�m� �{_Ϫ?���X����Pl5��	]�5���3Z-����Nw�)Q隶�ʂ������a���S�J�������S�O�����q"�Ӽr��"s8Y�Q�wK!�k��f��e���FR���L4�)᝔�)~��;�4���e7��^�8�dy��s����Tw�;�V���Ϊ�I����*T��b�b٦E�H9fV�֜��m�;�3a��L��KF�+�Ck�qI'��g`�ٯ��1:��a_��ҧ)�-�l�n\�������q�:��z���䘮ynO_��e�A~!�E�-�V�N���ɳ�N�)}���~(iJ�ߕs���ʚ�Uts�'�;�-e���x�}��+����C���e$�R��kXgT�r������0�@��L�V�5����|�^�Uv�!��~'�$3+��+���\���#�PQ��տ�q���;� �r	�ZNH�N�Ӂ�"�ͼNZ�m�֬b�b�B0�>�
�	���3�����v]�a�֬�)�B�x���<ǥ��'��]cH���e���.O�7�-p�����q?v�?�x\N��k�ZWľp���.�Jbל��S��F�� _��ί�����x�X�vr�W�/����S3�1׋	V)�lxk��5b��Q�bQ�Ka�x��ij��^�U�$\s�ݔ������W1��;.=��%�15��+q�G#���(����)���"2�^9�����Gyk���#Y��+�{��
9͊i�Z���Cw?�u�T�UU���Y�-��P�DV�ɉ�?�8��V���6�]p�2��l�N��!��k��~��r{�,.m�&�;��'C�n	(�M5|�K�[�2zi$�K8���j�5�?�a@������,�A�l��%�n�i����E�޴����p/c��`g�ܥ�y�v���_w�Q�z�������)QQ!1�=o�m�t'�^D�XQ�3LuLU��x� m$��ɺN�����0d�t�\2Qt-H�mo���'	fYи30��zc�r�j%��4�l>��ֆx-d&�������Se�S�&k��Ӄ(���.���AX�ְ�$馝�Rrx��������Y���y�&���Ɖ!]�%�H$�Cqm�	��xzy
��
��y��[a��5C�"���\��uCp�l��`d���AO� k�5 ]�K"+����w�3X���"�+{����ٿ���G�l~��Ri�[� Y	b�h��3��S��"<��~�થn���ޙǯ�������C��m�"��F��<u�����a49�;�V���g
��ʢ,]@���ĺ²t���%K/p���Sp�2/�"S
ywӕqm����#O�$��aw<����᝵�h������>� %f�V�v���Z�*���|j@U�ny���A��E�7���j�.��l�2�z��#���N��Ac3I��h\�V&=�\/	�_y������۳%��`Ő��%2���PJ�X����]�Q{H��w~�G��Ls	/4�ФЙ��͟t�D¼&m��](��q�0tx?�v���3��Dl�.t���O�c0Ձ'(�n�Lm�-m*�N��f��`�ra�N�6yP$��L­i�U�b�Ck6�]	�K��H\�s!����\�a[T�#��e����e�P��̽��9I����a��X����@�>nk���,�Ŋ`��M���Fx��+�ߋ�&v�'���N�f�4O��џ{���S��b��7pr݀י�����F2�T���~.��Y�KÃ���gڝ�W�R����;��|vfw�����y�B���D$x��1o�0�Ԇ��Ą �s����Pi����F��0�,w���
� �O�;��<Ҥ�Vr�9��#zbQ��x�K����m�Q3��Ï��C���s)g����w�Ʊ�1(��;�ɏq�4z�Q���gF?��\��8\��W�J�ރ��v�T�@"k>��X�m������[h@qE�ߊZjtn��#v��5�	E�s�2�
��Hۍ�+���<_�!�zJ�����*�
a�I��	n3 �.D`t�*�e�7`�!*�g�����cd�VF�eǬ{��!���տ�K�����VW�<f]|� i��~P:�o����m��Iu#��l�*���-(�*���"��(�b#��K��"��S"�D���A7w��é8qʌ��_ܓ|J���;l�n�����i�c&r1��߮)$��b��Ԙ2��,��ڪ0Iq%���%�f�3��'�J1�h��O�W��~U���
}�91 *�`�[*F�������w9�>z�`��pqe�N��?{��w�b䞢H�o�a�O��#�iڤ�$
���.G�N�xD(��w�n�Z�|p2W�&~\��6������`6w��F����%�&��C��,�j����2k_��#�ؙx����T��![�}�3�@�9����W�ˇ�����YK�R%��N�&~�˦��va��g��?��)f���^@��d{��g`t�޶r	<� @�P��/���4=��7��N�6�W'jqCH�6�Yq5L%^ш�!Z�j�.[��X��.�ʜHWDEd8i�Z���#�L:�%�>����O�]�3XuL.��w	a�%��j���+�#�+������j��&��P �	z�~V/;��Sm<ʩ�=�L��m�[E��ʹ҆πxdB����)���>zY����2�򎕔�b���Q2ȸ�HAG��U�o���J������I N��:GR,l�a^Q�I�{���_�Y��LO�`W���4�����_F�%'ݟ҇����+���z&')������ȟ�f���A�rB\M��F�l�%���'<Tƅ�����:^܍Y1%�۩��nm�UfZr��g>݊K����B����=����7_k��'��_.d�-��P�+4��^��N�q롟��*yC ��~N��4����Y{���T/P0G����
į���*R~��U�8�DX�8�:5 �p���ݕ_�����M������LSnRH�M�#��!�_��գ0�*,�bU��E�MW?�q�_�ˣ�װ����
 �������N�8z3nL|Is��!�*�p&�������]X��N��W�(u�P�\86 �X��7�5_[�N�FMb$�k^7�˿�lDr��0i2_�U����'��oY�v�T��(-);�5K�l�(K��-��C`��BF�v7�q�J���?/.-Mk��ӹ�NNYsOж�" m>�������ar��r�W��3N%��ffd��ϔ�g�&�����{���%q6����y�f�5t��*���.آ!�`\z���<#�X�	Ee���q�?�dxT$��@�I�$�G�X�	�6����Ε���_;��_���PȈ�t��*����@C_ki[l_e紽7��b�ʍP�b}=l*>"a�s��鋳�����%�}��� ����2�qM&+�%�c�E}��V{�a�b ��ߞ�m}0
�J���-�`�I���BȲ�V�8ǂ�Uh!��->~���Mh��IyfVZ�և,��6�/V!)	F��h�)��0k����Du;5߫bv�?�$�g���|˶�g���1�
s�Tݫ>�
�'�ǯ�J3kҠp��u�dp�_����?�w�	�W��fC "��]����FJ5h�9-h��$��e����}� �d����o*fP�+7%>���*~��yY��V�����g���!Ӡ�S�i^h�G����lcP�(P�<b�O�q.� ��rJ|�8����d�nB�G��(�K, ���Fe���	�%���<�4㝬V�O�lr~�H&�7��W'c�Y�b���PG�3ap�9�
���	��C���5��t�:�C�J��B(`��tnNL���u{q�SJJ�q����[���P� j^�h8uWj͢��а��*]����Wc���-<�3�gE<U���	��Ir�����f ����}�n�;��S��j���qv�/���y�DzI�+P���UY�_�z�������_�'���IS�f�ܬf$Lw\=�B�HxWr�O����_���N����VM���:X4��'���{��CQ+��)�/3��O��V��,�L��gP�����;N)��EtU&���F�߶YU�E�Bt.Z�͞!h�ݮt���	v�H<�$ul:�?�Z�+�ꂴ]���o"�p�y�W��5l�%�{�U!b�洀�$�rd�deü,˝�g��i�0G�$z���bi�~`��
#>A�Q9?�5������4�	L�Q�f1J{�乐{�r g~��=��o����׌���UЪ�����`�}�B���h�#�6�		R`d���AW�n�qYW֨6p�1~� q���#�ژ�����!��܍.6��P��125�&����9]k�ɛG���#qJ�k���|M���#*tB� ������}!�'�n�lނ/��pY�HD���sXa��gӓ�� n�Z5�b7۫�-aRf��.�\�:��>����Q}���=���Օ��/��)�
r�ٌ��د�܁v�	�t��X��BlB�������=�;�\�"�t0<(x�i���i��]��~*h��g���� ��3H�|�~�ʫI��\�RA.�5�#���M��A�I�pw�,K+ej ��eϿ�5;��XVD�+�6�!/֓�5�(IFJx��Za��sp�̢���83��G 䖩b�B~��ũ�De[Mx{�̞>�BQ�(Ms�t�M4k�
����r̻g���LK�ha7��i�)dؙ������ ���(Vg���q;�wG'�}�q͌��0 �Ѯ�|���N(,pmzm �1���xq,�Jox�����hb$��3r�|�-�o`�������$GH�{$_sp�q�=,ّ��JmA,��R)*��V�X�g�o<�'�$�v��yP��eP?Q� D2�'R��'4��2&�S�16���-5Bp��t8ֽV��sYHO���Ɋ�f�	�ON��D��_j�ϑ�� ��L7��@�hD�)F�s�V��eS�������~��m����c�J)��s;��_�ItԜ;�X����"5|�.��\��U��h�u�.1�Q7,�X���A��D�17���"�^�&D&�on��C�'�KY�A����ޕ��ԎS7I��h���r��}/����ވ8����l�q����vX���R���2&!����,i�KO�=LBM�ѥG��m�n�XW��& �UΙ/`�PV2K��%bս�r���䧘���_�(=P���[lYr>�`�Z�"�tĥ�����>�)38�JBIiM��W���M90'=]���9�����'��ͧ_M��,�[)��u5"�F��C��^Y�Q�?�̷-�vBqt^�����m	� 6Bt]�c]��a��� �Ȇ�,l��/�}���V3:�t?�\��EA����{0������&��䉄\�X�ϓ�)�*J;�+�+3�D�Hd�����5���J��X4�S�w�r8����[��a3I�b�d��d���Qn��sB����d����j���>�p>��:��4�'_������B�^���겄p�dD&�!���l:��J��X��d�-o�!b�<��v(�W�XO�7[�3Y��B�y0����z0k)ȷ+j�q�h�M����Ň��]��q��o]�{(ݩ�a3�%�����|A(��
�[&�Ir��w?�k�%�� ~(�ڽB�h��R�%�|�����6hV�����WƪP�}P��i�X��Ċr�n��F�VQ��Y��EZ�k9�t7q�)(��yy��x��@��;G�FT�ⓨ�'�ڌ+D�`w;��HK.<|�rN?k����*���=d9�a����TīK����r!��:t�����+��� �-�`�Y�E�C�q���{J"l0�6����X���P��e%v�Zױ��=&]���E��T:�E*��28�\�	C�o�BioQ���A��6��S�EA@1 ղidDMVP��vc�����u6[b�M�L��D{����mNw�%��0S������(��)��!1,]�z�h��,�)P��XH�ؒ��@Ƚϓ�O������s���p�����o!�~��[C	ᭀ9�U�|q��{��A
Ld~�x&��I�o����$�P�߲ɂ���C���w�CD��t��ݼ�5�y��{������]Ca�~T�bc��Aq`�֌�6u�����5{O$���[�)QU n`\�d�;��M��ha�� \�rX��a^\ΐ�@W����׫e��Jp����	�U�.i��W�(��ŵ0	�݀]��V��LbҘ!'(*_0����������na�'��0i;r���-MZ�D,FΟ�����S�Ε4hR�'H��?C[�\�����}]�]g�x,�`��21r@@�����y����$i������z�9@���xM�go� �bx�(Vs�t�f��L�C�pA���\���?f��  �2�?�f�^�3���{4(�~ |��Թ�[Vq������V��IS�\���"�J��}��I���hz��q,E��3J;.��X��C�� ���]�lÆDu��������-V!~�OmɏW�,����E������$����|@��	����\ҿ7e����М�V�m��2�d%�f��J1����M���	���7�U�6�L�� ��<����:���#��juA{<�,G#ZV�	�)�є��Y�2���~�C�E�㮗�з�$�RROX��kAR�����C����F\�Tst��v]�z�xڥN��B��*t�D�/�"�0)^ߑM�������A�:����-$�sZ%1���.b`�>��;()o�!��@�rш��Z�]e��e�-[A�a�����*�V� ��m��H����;\�����}�R�O�F�ڹ�s�U��������b:���a��|�-��V��Y<��V�=�H@b���3o��SQ���\Մ</4�U�9�L��Q:�6L�RgU���8�D������֣��K����G�m���m:�&�2a���.J��J׬L�ȑo���-ѵ�YYgԂ��������M�Aj��޾�7����<,�����lJ6)?�@��E���8�9V8����:��h��ĭ�T�/}�$�)����!����A��[���3$���@�\|J�1�.;�Tjt.�#R�퍒̈́����P�h�PB=�W�(���j�U��C��y����T�����EE&ԋU��Жpʝ�p��-K���a����~�[O��������@�^7?���:\pC����f��3�3QO/wG�(:��T�L�2���gy�"�R�^�7���B�zF�5C��7����b8�_���3����T���e�����\[ؕȇ�O�曺�'A��P>޻��8��T�R��7SY 3Z7x����3{�
n2R���^_�e�;+�iܗr~"I�,juȎ��Q�y�GJ	-���ȳ�-�IR�v��&{z?Fq��Q�_�w$�$~�n���D٪�
������Y\�]	�j	´��Ѓ<�=�F5x���<�z����J�J��-�1n��[I�Ct���rו�����N%dLʗdv�0��i ~�B��j7KXѵE?F������/"��/@,(�O&�n �e$D��0�x�n�	�_���u�[Z��/�B_g�%g�0���:��4����ʀБ���[��g��:cr�C*�嘖 !N*;�='�i�瓮3d	�L&��ei�O
5֧5,f����b�p�#3*ܚ�)p!�����W���MA���8�*��3￠J�Vvu����`�i��{�� �_��܅CP)���!��[�vUJ �=���a��)�7� ^U_K����17��_>rQ7WP�twT��!�2�YF&��Q~߄������'���f�,ʲ��2�R�;�ގ
����sc��:�$' �ȋ�h��gV%1Z�Ê�������od+��Q���S���҆�~ ���Gs�>�)8��b�U-�]���X��'/��Ù�x�߼��M�(?_C����q��d@���7�Ԗ�]����*k�K��{.<�����`r�8c��KY]��i3�-���i��!=�(g�c�NGbӠ��oՕvĔtZC����:/d��='�C���ʪi*WE��<V�Ta�Z��^�u��> �(x!( S�d!l��)BS�~88M������rG	7���@����O���w9�?�M�����\��X5p��$t��]U'���gC4پysF�o���gI��'gz���1�Vf��@�MIRZ��/�*��⾌F� �T_��ɵ�?��q�xƪ Q��e�k���8������9(��J>�q�IsA5SK�YhS�s9�������T?b�Y?!��I�I��ً��fLRo�j��$ b$n~@�<L�

������WYg�l������T�Ͱ�4�dك��qi�u���O;C�X����*s�ɋK�&�i�&�����j��8b#�CB���r�,�C2z,q��@�R��Xq�3$��ӈ�����S
�~�^ARxh2@��D��|y����_#W��b� #�J2�
�8AϺ��%@<5����3����8/ay�F�8#q�b�s4����t���8�r��h��0<�<o1Y�3T2G�
���J!�(c�[��f�¨�^��s��wT�y9�����E߁��LK��ݰ��?���*��v�d!�*L��]�Z4�rb)l�}�,�b��N_��j�Gs�&�!]lZ3����i`!
�*7t����Z���ED�ρ�e��"Ճo�h����Y2B�Y�o�_��,��b��g�j�Gi��S�[P& �aŦ=�zLx�
 ���Vu�ԁ���T�&���Z"�t8U~8�z��_|p�
K��߅K�9a:��f����	�鎏
���$�����$�a���A�RD@�c�ɥ��c�U
��ތ��GцDy)Dw0lv��M�XC�m�s6��c�lS�����3��
r����=��|յ-�tW���%l��|����3��D���Qe��F�#d +j�˃��|���:�`� ��q�B=0;=>кR��A��dC2m�_)9Ǒ\���k*�3�%���B�0�p�hŪ:b�R!�+�X�Y��i
CW��Z$4����*��O�*����`\F��\��1ׄ��	?K�3~&oYu�컻.����e�?�P1�D�C�jL�;fw1r~uF�#�!�t]�?�$��B:�`A���Н��$7p��O�O����@Y���pj��D�'�}�3p���h��_��v	�.��]���E������)1E����P��y6�?�6&A��'od�YⅫi�+���쭅�+K�� ��[g�!r0���G�ջ�~k�9y����.uƜ�}�v�Ư?�	�u��H|y��,=E�>�"%(���"��<#�,N�'7�X�g��cb�m6H��2��W�����r���[�����^�88�����-ډ	�����v��Lk�
D���,��������#�S�[B>�8ֳ���>����x1l����/��X��p|����F��$����#�3��jE��)ǈG'\(�(�U��t��wXÊ���OC��3-�# ��K�l.��2�6}oŰ���9`�����՞_R�rR����:�p,�$��T�E�/?�m]n�ʤ��/8 e�����dE�?��8�L��Ae�8 {PϪb���c�퍪�����c�����߀��ؘ���� ؇6�i�D}�sC ��$_0���Jc�!�'�M����������w2��|l��Nu�-yLy�X��p�4�ev��
/�a������uUJ����Qc�c�Z�J��q���}��w��S.g�A�����]���cd>�n&F}I�Hy����&����XU����l����J�үr��x������Q/��ٵg�[i�7R,��at�W��#L<���^�}[`_�o��No�w�`�3S�n)�{�T�9����*��V����-���D���e��H���>x�>�a�ie���R��y�ki��)!>ԔYmp��}$�𞅂xȸmC����}!�G���$9�MliՇ���f����\a.S��%����E��g�Kғ �i�+�u��%۶�����K��N|X���M���bR����Q1�lq�	=)�^�nS�X�)$�(�s�k�0�h���/�;�]���'�sȀ��Qw,�uPM�nBF�M����s��W�5���5>��>�V@���D�׳j�+�䀌F�r�T	�|�^���m�����B����N����]��v4��)��
x�8L�ԁ��=�V���@���dF�O	�#u�-.��i����B�zM�m��V�'<�_$�¶8P�F���$��Eq�~;��bB-��´���p��I�)V��4��Q�S#ވ�np�m��� �P��`Q�>82LL�A�~����p���Aj�e��]�X�n�>��ك���T=[�92.KH�v�0R�U�����7���O��EL����[L�����A{��1�o�J�����<b/�Ł�Ƈ����1��I�RFKv���wVlYԑ����|���_�#8������ms��p�����\\��V�EYwl.϶�Qx��׳��b�K�PO��2�TK��?;o�m��c
�A���j-s��~Y�'��5\���R��~��(�S��hX�B��3�,��<�p�H��e�h?�Em<����ה�|۵����𸽐��A���E5�Tq�R��M�?3����&D_e�K����w�_�����}�a�m�k�jy�$3c1���Q�X�޽���ӄ"����YAM���BY
����O�jb��pś!�9�F^�M-��7Ȼl���q�+�^N����A����vs�^_4ω��J���"�L:������O[�O���ɹ���gBG���.�P�� ��H�Xr�މ�un�6��[Ed/�{�&K�����tb�B�����A��C{/Y�H}/�s��Ӈ.ە�:���� B������v�Co*�Lc�cO�δ\aIֱn���m��vtR��v�c$d4�8͛���P���I'ܨ�۵a}�z�T
��0V׃�V�����{Т|�Yr�W��h)�Ї�ʜ9FL.��R[��N�n%��x����X��y�&:p��p�� *��z�F=j�(?���[(��q���4�����_���4�+�\�7��0{@Φ9ѯCk�YH��e~��_Էq�T�4�i�5�` R�K<�.M�;Z�ͳ�/�W�+9 3����	�5�\PE������f;����l��]�j��.l�(�l�\ߪ��d����oO�ũ"�Vd����1�I!�_�P��#*?�N؝{%Td����v%d�?���I�x���;DV��߰�)C_S�g�oj�}�+gp���\�C�9k���X�p�y�.`:���J}A���N�"�r�^،�i��F�}6d�
u�"w�)�/3�����wT'�Iv=�,�����+���F�]t�1���7�ԑ�i&E󥛫URv��䏏H�wn�3ת��K�s�,b�Q���س�qpDI�р��l-R!� \O��nY/I]�I��x;�I�|����8$г��ᮟ��ǌ����^\��Խەqz:!�yA��$~M������#+`�''�S4�"��qS�ij��L��T8�f<g���>
��)�ݗo��Q$�!�0fk#���«���Da��-�>e�<�%�z�o�QS�ۿ|B�_.��{��J����3��'�'Ae,��}�UoaFY�����=x}�Svya��|�kx�\��j����^�of�˹��)R���ql�3E�b~T��wԏ�?o,��>��m9��8���o�A`��l30?��yz��h��;��o���᧮cxE����RD����pm`9a��M�[x1�n=/ަM<6T�\���ӎ1?b�	�[��/<�Ă�=������y1$�M��"D#ST����fD1����ʜD�_��o��E���	-��_;�S��3�+e�P��*8X2������=,��9k� ��ڠ�c����'��l�g�vW��wW�%�ρ��PJYR��WN$��x�����\|UuMT���=�;��RȲ�X�����e�'���i�Θ�w��`̾��~t�)��?�20%�&j|��w��W�U��lo��E�C���^>9#��T���W��W�L��3^�����nG�EF���ĄB�8��D'�j$\��JXV��RA���s��,��:'ѸKd(��0���Ǉw
��5O�im�����Rs�_@����v��V����p��˱x���{h��MT�zߕ-�q����62���h˦FE5�:f��`^���^�_5߹�*�X��W&�C����ޞ;焐�J�.��oE����G̀�WOx�ǉ��^���ƽ��wDY�#'��#H<fҷ��7�[�)�G�9Y_�e6�
�.�[��������_G�o�X��r��̀D@D�c�}#x�S0�'
�:1%~E��Μp��S����cr�)�R�Kro�x$��oVv�/�R��2�݂Ʊ�K�S�q7t荁\���F���4'O2������d&�F����F��_��=_ˮ�3�#��u�c�^6�һ�a`�0.z6j7h���u���-K�"�k�-�ǖt*��Gn�Z���듩�ʐZ�80��%�1b�ڌ56�����"�ZuqZ�J*񖷔VrE.��a�(fg�,>a���_�˗�N �h}�j��8�a��w�D낁v����﨏��x]b ���B�p BZ��Si]�y�k��P�;���Ujbw���3���h���Â�pIs8�
�����Y�l�Z#o�w����H���F*����rޚL�g��\m|��cs���F�6Qr�hLj���m�F�k�[0l��u�2D���Rx�+tƔ3β��܆��OU�.K���oDM��-G����.��~�@��$��^I6��
u�"�脷s s��L�]����Q|�������sD;��i��D�i}nD��˯����;�Y~t^��̓��.3�* 	8�棽�=�z��|<X�N�m��M��1�E�o�/��}t���v��i8mE'�Id=it��g��oq� ��K&�ș�"�92h�ѥ����8���fu��Ȱ�lʵ��W�,��`U%ߞ���T�0ĉ>.J>h��8��{��"~
�9�,N���Cay'���|xo�)�%�a���\m��uuY����_��?[�9��ƛ�y��%�ez��cՃ=�Oڜ����F�2��OP	kIB�TpC?h�qS�JpG��|���!²1ډ���>�@��s�o�@��o{]Q������c^5�Z�#&�E�҃��g��*tb� �A��[��<��4�W����@�8ݤ1f�(iHF��ڟ�$��H�;��?Q�퐥�֫����`݌J9��}g�� �ќV�FDv�$([gXy�캹 q�j�{ŜK��Tj>�{p�-z��N��HB�F�@��U��)��>��~G�wf���E\�W��Le5��6����cڴJ������g��,)I�D��a��z������\x��!;I%$3i��/i�!�Ѩ����V�]������m � 48v��(L{/B����~eeߺymx���p���N%6l⻳�W����uB(7��)����'Y`RwZ� �t:,O���5�i�](��Ή�`IP�!gT9��qI@\j�3��)`~��Q��?6��۵&�rj� �i�0=L	��>��w/�ʑWdS�z˟�՝�W�߾��;��Q��\CՀ��v�U���G�S[�&0���X�;� ���cJ)�\������{/��T0���7V��e��,Nn�b�uޠ��{����м�SV,���70��"�$;���y����Χe�4��s8(؜;���5(;�����z�5�Ԣ�D�k�����/�rCQ��[_~��f��KHRV��?pW�9
���{�tݿ���᤟��3?ۄ���e:�G�%,��e(8!�� %c�Z�o0>/���Y����U�WO0���.g�o@�qʣT8?�ҧė��%�b&���rQ�U(�Gtܭ{����斗l?7�zOl�<!�����v�ė�z���\����и�l���#�R�]`k:m�&��h�`sب��&�҃��"���(���$-��Vϟ'AC@�A'�������Rs1:/����Na6vh����N�q��Xn"��t,Zph�ě�H��Q'N��4%�}Y���<��k�!}�[*��D�xg8>����r���(�=�k���i��L���^6��lE6 ,5�7�? ��*�QQ��-^�9�vh��5��{�50�51��!D�����EbC�C�$�.���
7�FJL�0i,�C��7�'ͥ*��8�ř�+q0ZJ�G����fiP䡀O8�w�/�F�=����!��#�Um�Bɶj����i�Nl��wD�
I�����a��'��j��fHy�/o+8����W#�;Q�������Bc�@��[��B`J}F�wp(��
&�߼+��@�� O�0����,���轐�7&�u�����0OC�L�^R]�hM��N�30�2�5D������֓_���\�Md�J�uj,�e8uVso�7�4Eq!콦��k���v����_�[�}�n=�����?!}�o���*��/���t��d.>%c��6���e�]:%����z���ņ,�r6].�֥<\�]� D/\�6�9����0�>o8��,�f�/gK�r���:�k��$������G��̣lp�){��8l���鴢��X�ޒ~<�'/!ГG���=�Z�a1v���`Z��n�{#�� ��;kNpM=�`&�9�Jx�e�Y��,�恈6fD�E}�%�'��̙�=���ʝ�\��ɃN��A@Wi�_F������g�6ݶc�c8j��(���)���dI��)�<G��M����C�kZ�!�2!-	��[>���l\�A$�	A���N�rK��p?��SDf�W�n�SV��T�M"2���| @k~ӭhK��}ӑ���
EU7��M.�\f�~'#>�R���EH�B�~��FبP��i��ʫ�As�j<=0�XX���d|~��nv���jp|��'䑙d������5q�_ov��T�
b�� �}�
�"��h�c�<u�O\��uy��+��X��^5l��%=Pv��F���!�ekd�\��;��|(V��1q%P��HmBd��HzԺ����k[ك9.�P�J�m����@K:oB��)�`ɠ�L���ap,�L�=�3�ɹ���z�J�u?mf�!=�OH��<���2�<��l�Ɔ#�d�-��%n$T"�p���O,��S궭�T�Ψ��[�Y�,G�Ѹ���N!�����6����/����������I���үJx��!��Nߔ�N�4�;(M� �]��ㄾ�ʊ�B��.�i�'�'���BO�y�[w�5��(�
��&�0u*��ZZ@�,��B���*���N��w�H�"W9~#Xo���&��*F�L�J{�LC�gJ*�<��3�����������1&�������YDKrT�� �i]:�.T�[�� ���3���R4=Km��x������1���Xyq�HW�����yh�+��]ܒ�H`�NE)�2�&�TM��`�}�Y0�$�lu/&��m�A������K�-u����H
��/��j��rjc?�]���!�J��W���-J��jArA���}�v�X�R�S��s� ������J�%�J+�ʘ
ɂi<\Y啲�ʏa�� �4���Jz�WåM�o�9\�����Bc��1O(��h���i��p�I�0Y�������bAJqߣ�]*��L��ӝ�����U=	�_7�)��}mt'�����n@�TYH��#p�F4�><��8�j��|�-p{�A;��uQlC�'�]�=`c��LIl
��e��9B���� p�_M��h���"���AWq���H_(A
�F(e�o�%/j
R�b
���_d��u��VeД�����v�JSCw�Cg����e�c~��ț���a7Gz�<�U��&�/��"�.�s1�x��!������ܘV康�|�D��hϹ�,@�ք[�ݝ�������2���Z�4`��7�|���N�ͅ�ضE�r��2+������˦qV 6r����+��q(��*��۳�;K�y�L�4����l'�w W��N�,��%ӌ��+�y��FN�ȴ�Ch�ߧ,L�p����ErAY_���@��$�P��<A@����z��0�����0�n�}���4Q�ڭ���z�u:������V`�����g|�����Z�rB��S�g朾�z���w��
�:�&Vu������.�5��={��0�=>a7�=��B�P�^�"`C�-	�&o��4����o�N҅ZY�A���,B���ܱ�+�"8��?U�9-LX�q�*�1���z�z2ɜ>��������\��]��l��3��}��>��������c��$E�J�/�����"�ml*U�!����揅s�4�m�9C�ળ�[�&�⡈���C}O�&��hA�ס7�$��`�KwW���� �C�M���T���/Ӕ�S?�9W�M�I���{<�����k��K�D@���N<��,���HpQT3R�WJ�ƞ(	���J�����@9*���~�d�s����es)�jvF!,6��Kӄ{u����Y�u�����j���1P톨RR�Einnq�/�U5����M�{#6p#F�������K�׹�<Gt�I�Y���b ݋��<d���n�т�HT�:�ص��ìT�1�t��2>r�0:�{����x�y�*�a�:����'���]���^A�3����ɣܴ�)�R�*TU���/�:��d��^ٹ������~�0bv�k�S։Վ�6�B���$����Ȍ1�FP �1O�]mصԆ��������r�z5�������D�;O,<`&��w[=�@[=�JbH�q�4QN>���b�
��j�ɢr��B��;�?܆�pr�ؙl��k3����(���Ю �����9;Z���׏N*F��!�E�t%��~%�S�`�YVq!e�?��A�� �T�Bq%��'��Gb�?s/6h]4������x;�Ra?]G\��7�:ܝWBf�a�M�$��`)v�oe"�8���,�+�Qs�$'ޙ|?�p����Hۆ;ೱ�{��ا�:r�̅�ŷ����M�	�W�r�1[����)Q��I���FTY���;�7�F o\�5�T�:����yu�=2 N���\��[^� b#�kó6o�� ��$Mv��5�rV)�)l_���i;��� nT�3�<��AK��L��-��V�r��Mf���ԑ�Sy���aD�7��A��� \֓�3oH�8LuN�L�I�I{i�������O�4��r�&��G�z�[3�.Ũ9J,��{3$�E��\��#";�Wk�YY��FoSt#R߶�VV��y0]���d~fg~qaj����Y����m:&����ʖZ��cfX���8x��1�^q;��@�e?�-8�*]I��]m���y��;ո�+�-&<S�BPn~��:)����&f�jD�'rr]W���nN�Y�	���{��Ԭj{y�.{&7KC֪
We(DJM�Ә�N�I���Ɖ�8�r~`'��Ux�����ı��x�j���W�l���h�;��*���G��q�6 �$e�g��J��`��WѴ�:��Ȧ�yQm��S���*L��d���t:��_��k�g8ۜj�e�KU��2�5��!�{�j�k�S�5��0G�m�Ѡ.������RQ=^��ͤ�>\xCoQ)d(}e���|S��GD�ڎ`;M�DY�MD��P�0qv���i�I��X��3 ���k8���R��M����4x�hdjm���V["��;@05x���n齎pm����k�JQ>�E�B�n��Z���[��vDeh�s	�}����׺O�I���ib:�
$�o���j��V9��h���z�*�$ĥB�i��z礕�f���bD��@8��
D�d���C�'e˸.z�I A��0-��D�"�q�7�]�� R��)���m�q��W�Ӝ�D��&���`��0�FV#'6������>�L�.0c����$�I�ɉ����?��K+�H�<3�@8��$���R����J��,�;
CNt:�be+R+�$�)'u ��Pl�Hѥ76UV2���g4���a�?�<������j=����i>3�D�ܩ+�%?���$]Jf]G'j�6�UC�.ɖm�&El�t�Xs����Np��Qs�>;o_�t��z�.M�Y5��Y�h}�Ҡ�ԠW����Ϳe���r���n	S�3��Yb�������-<^�c3�y��A��Kʄ��)t�Qp2|(�7t�G�e����kf,M��b�0����"���#�.����rE�dc�0��ud[E� ?ȱz:&��CFo����"|0�U~�9'��V�_ڴڥ:K/!�j�ؗ����V��M=�͸YoR��z{i#�J蝘�a[�8�F�Π�t䄤}*�2�п�]������	�7�cH;Ƒ<�%b�� � �䂝s�Ȳr�W��$y�p}��5���.~!��z�o�e�����ݢI>����+�"?��yf�4I_��Uf�
���n�^J�؇�y�*q�Z���h$����?���^�^�����|u�|�iX@NT|
�������85���A�=���A��ض�U�l�0sW���5�0��
Sa6�Ȇ{�h��N^�0䜞\*�Q��M����������M�7b��{ Zְ�Xm�~��V��y�w=!xT'��{��L����l�,�ɐ�񸛳=�tȐ�We)jd+E�P�\�|�x8�����u�Ԟ�k����{�|�';�E�sYG{�9cЮ��wD��bh%����U�p��8SF�6�>�p�ھy��y�ְ��ځ�!�}Ѳ[�DUWN�+�� �H�������QRa{� ��R�,�%A]�[�tՐ6Hz�Z)��t�KI,U���RD�x����0-�|p�;?�P�7���oE���'�T��CS���A����,�NMf�������T����$���d�R����M�9䎪gY��P.�C�^s2�������l۵���J0%�e�O�+��� ��V\�v���S�Gd7�l��Ͱ$�l�o��)��U�/y��d$�W����=����]�|����fd��\��a�v)�:"�@�����1�F��Ř�QYo^6$��1�0��@R8Itm�0m¾�{�WEz�?��U%�Px��� ��\%Mz� h���
��l����� \)���Ÿ6��;!4{B`l���E�JN�јU�./�n��n�`��	�`6C���:
��28rHXҡ���ɗ*�!�d8�҅)�L�r�t��	�'U�ӆ��u*Ծl���L��[2�^�y�[ڦs_s��x�L��Ĕ_��~��e���%�l<��vIQ����@ߛU�Q�Aiҿ�g�m6�TM�qF��sVF���Gi������)�����oK݇�TA��/,��F���*��lu&>\���{�0�Y�bgW�����i�h�3���9���Z�� Tm>5x4������!$�jȑj�����������ƙ�H�3�T�.�`��qr�ڛ���R-�$�+�a������o΄���+%�ǣ�
fW���1n�w�Dh��+`�@(�֝���lA��y����H�sI��^��I��3��r��Jݟj��.��ZsЮ��k�}al��Zq��E��Z"B��ED�|̉8!���)?$���4T^3��u�~�d0�Y���PAa����0�Y+��w�A�Xc˔��}��ߒlJҊ�3��w��MU�ۑ��ˤ�u4��M���!f��"����D��d���Dx�r�`jw�D�Xp�'�����&��O���ڳ}���G�d�;o-�A��T�5��e2~w�70֯:������ђ��T��ʆdg����m��'MC�=[�p5�<93b=�}x��p�L��
Y��Օie�+'!�L��^}��x����]��;�Т���`�vAX�I���\�A,�t�@��_�,��� �OԠi2ї�\�������R��X��ot�ٽ�S@�,�϶�i�[�n>HJ�7����g��y��E!aOH�{��ʕ�燑�N��SA�x�-���X�����mV%0BŴ�B�f�[-u�\a��t*ӎ ��<��!�E�[��:aҴ�)%����Z�&�?X	���GT�%� S�v(A�ͮ3���׽k̟�뜑r��E�0%��w<��p�(�gcH|�/��{:�o��H����V����S�X�6���fb���p"gw�u��X�\�ۚ�j~Z�J����<�$��|w���
���Cx7M�9=��j���+���nn��w��\��T��ѻ4f��h�'^��N.`�5�.��o�8����-��a�X��k�N�J��!'��+�S�8���щɀc��A��q`iԠ [��������E��'��Q�1~T҅��`��8v����H�D<J{�L�;���`�|t2A/;�Vt�[f˱ph3�cw)Z�mnHk��j��9�ӨU��n�n��
�>�)|0^"�tl|ʉ�
'�m��Z����U�������9��̳.�[f^�eN^��T�ԫw4�y��q�m%|8Ѕ���q�ۑ��|�8pN�q����h jo ��� 	�+��(s�H&!�_����;FP&�RF��n���+�C�^�Lzc����M�L�"���^.*�PN�;��9({��AO���Z�� ��Ä>t-���÷�F�����W<y�pQ��]�EA�Ԧ=I~���)���Æ���:�g��;�CV��O�7�N<G�	B��0���[��W<��I���}o��>b�g�`;��� j_{�&��6��i��9ӷ�����L�3e1���!�C�jOe�
X!��s�p������s�5c�-�]Z���quKN0b����e����^��} d���d[t��G�-+�O�qy�gTwdx)����xS�ϯ���%
s%��x���a̋�LͲ��������>��R�(i�n�@��f׬,P+�B��+�+�̛�S�z�rtW.x�lJ��٧��먆�KEV�6�N��I]}j�2��Gh������<�\v�X�J�[ʽ�\j�O�D���@�ג�i4���k�J;�P³�2�$;*|�x����b[ Z�i�ɻW�x�]\��tj���+��|T�vmkX�aH#Wc<��&""s������R�w2�����Y?��YA�J�H��.�}B��w�=��_hgAq13@�/#��r�v��n����^�"��y[��ܭӫ۩#@��R9���qr���S�rҦ��vT�n���������H���[�X��
>�a
�uEȬ�c��5Kk���)k�b����p.ߍ�� 3��g�-�h���	���G`u�~�+86�t,�$*,#��~�N^��7�.$I�8e���3~�١�RJ��ѯW���V`�V���0��j��vv�j[���=h=�����_���14�Ԋ����;ID��py�����%Gz'פ��0uL\*��-�?�(̦��H^�۾3��NF�(���������ʗ��s6���X�[ٔC���u�u���T}O��7��:��4*��	s�ۇ6�vy8:+�Ѭ}��0
�/Gv�:�?�d����|���KM5"�߹��F�ƾT,��z)-�B2P~�(��S2r����L�������Lc����Y�V�6~s���3X�S�����gG�վ�CK��b�y?;���
��ϴ�a8U�Q�+-1����%1�}�;�M��e~�^������^v)���"̴>�o��&��o���p��j�U酖�[��GCef'��m\m9
��a���Q���Y�`:�>�$'z�uO���U{�q��~nn��u�v�EE-^��:\��i�g(Ӗ�����,��ѐ�;���
�}�����]m��=a6Mek�fDz��f�S�V���`�Ki�bH%}��Dq�[�!=�6��@�5��Q#	����Vʮ�3��1r-������9x�,[1��Ա�n������T�}}ov�`D���b>�Oy�������EE�کR���[�&[n��_m��<�T�J��0Y�ߡ��Ɨ�ܩyK�Α[&k���w�5B
Q��j~&k�6�[�F8RQ��.���@@Hݡ�M;{!������fѩ�%�t��ncL؃�a�`8��(#����*'v���'r�-"@i���쬹���µ8��12u���[����~O�����{;V�ĉ���\G`�!3/�u?�m�����7�9P�6��K0�G����L�LU\��9�0*cȆ�����.��h1�
~Y��\�ع�A�
A*!+/�2�j~���k]�k`�Hh�j����B�ťM��w�5�
�1ί��X�4ݢ�`rx�ϧ���\�!R1�8��1ok�P��2�(jH�p�v8�W�N�3&����0�5��!y�(�����'�p��|��Üp��`������5Ї��c�>����)0��T�&�o4��Ȝ�Lz�D�ݞާ��HY�`�;:�O#����]3�F���!F�^��Tψ��{� ����}no$[:ZJ�����B%i;Ǎ����p��Y�E�3R�]x�ڃ�x呉E�d	"����2N�!c�����{�u"��=���) i6�0�����?�����,7������;wA��'Gn�$�V㫽���̜��V{7L��ȗ]3;H�Z��_��M�Y��L�kN�x��Q���,to�P�k!�S�_ߣ��SJ�!�My��߶v�o��0j�wsu� �¯s�k#�RA/7�Z^ �����-������>�
��r�ù߃9����^���L9L�P)'���w3��f�]�r���m�)�Q��jͦ�q"(��zC�e�P_�y�l��O`�J[��3p�M=�q�G���t�u�d�6疍.�R��<	��pi����+�H�`�������Q`+�ÇF	�
�<h������T|��s�ij3� eN��a76?�ӴXrH;�M}@�:�����e=Ě�AY�xշ��d�q�~�O�ɤ�g�8�p��4�u�tǕھ4w�w���Z|׎/ӡ2
J�>8B��R	�����ݻ�V0�N1��{��jʅ�8>/�����+�7i�I<k�d�n�V�jD�D*�t��oN�й*v�u'������V�\ϳ@BU6�|;n8�N�t���W���)��*b��DY���7�݄ӷCtH��v��F�0�Tl���;M)�����J�����W�T}��h��q��C�Jџ�OҢ�'� �7��֪�53ފ���٩9�W��M�6K�e�/��E��K��Ъs���۹�P��Z��ۑ����{�h]��X,aX���
��g��%�1�M�OI\��E�f�5^�<�{�f��X���\s��˾_��	��'�%��A�sK�Oa�ì�����p(~�Gr�Vm��˝a�³k�$,Pt�x�Q�4��UW�
Ei[�è��t���cf��!ك0�|)(g$`�0"7�Y��3,�z;�?ZM���3��w��A\��`�iθ|�:O�����52��d�Y��*�ڌ��"
�}e�n�G�Zx���%=y}��-_'R���i@3�_��6�[��Tԩ�3�9��#�Id����a5MPTAS����QqLk�PG�8_��U��V�|ui~��̣���/�s��+���p�`�YP�5f�7�3{�$a���&'�d�9B��+o)[�A#C�����;vy�na�;���ʹu��6�8I��8�X�^�<D��ߐLL�	��e��=f�2>5��hm/���X?�O�YT ��0����x/�WƔA-�Qw�7V��ۃF�@hi�Q���wL���0�9)����]*��91-��C���!8��Qw}�]���� ��N0������\U�D��ߵG��5����/�u��l�T��� �>����Vf끃�j�JNx�+I~�>���)��sf"r��$�Kk+�@)��]0-Dc�!C��>W��si�����Sj���x�i�Jo1.�}������N�!"�B���;XĚ'@���H@�B���m�Q�x1lE_b@����r��z���%qR��O
J�۲�����þs��?��U��{̈K�7�&�a��g��,;\MM���F����g���Z��8oǞam���{�i��I,3L�qT��Ԧ*\��^�y�kic�_��&��W� ��AȐ��52��Ү%!4��N\��t�Z�0�f���GЪg'v%;r��h�NOe�3Ŵ��۟Kq��ѥߊG�*a�R��z�����s��z��ə=��}�4�"݅ `e\���5������nS�1*|	"�}�T�b� �!@z|�jH U���� _�WK�nQz1-�F���d���}�D��P���'����`(@#�(��Fo��RF�����(�İ:<��-n���,��\�i?�_�w��J����G�w���M�p�:���<p�iR�Ȱ�XI<D���'�N��E!>{�4���~��'��1;��:8�ې�$5�A�QS�*1�2_�:��~bf������`��;�ClA�[��ԩ�i�F7Q��V�`�Ͻ�K����g_�r&|q��2�_G�R�Gv]<5"ф)/6�	�ƾ@^�H�6�jS>B#��{��C�#8��r��7�*�@���z~��C��W�(�!R�d��1k�
�U��i-O><;������W�~��H���QW��Y6�0�me0��]Hh:j�cv%z6s:*(T�� "PK��Z2�Hn�ͥy��F�5\��-�@u^�/^��{����b�k,ܩ���S��@a���1��t]�n�UF�a	�?��!,������X�m�H�9�,p�6�&��}Ϟ�����4WD]�@K,��Ｓ �J�`d������%C��u�U9�}$?��A��4�!>�:���nh�@�_�b�I���[f���-�e���!"t���/��س;�L����k�Ev;'�j������$!�Ze�w[h�j@G%K%����	=���6�Sںh�}2 ���؍����s�o�� �;�F.E��ԠhFG@�QxO�|X3H.��ňj�G�����WÆ������:�]���S�_�D�v�x��>V�2��d�12JQK�s/<= �>����b��Ua?����N� �&}��./���9���d�=�Պ���%�jd���9AԚ1��\?�ՊյdW����`������M�3�ݲ��h�/bЂ�>CkVRR��~��o�0GLJ�V�Eh��]_tO�"���������}�6"�pF�Q��W�Ba����{�߻u	��ܸ�3m�2B	𽲬g��oR����Uj?3�t�M��T�����v�܊��S�O�#�P:��i�f")^��(Z�YWi��y�i���f�l�aA�W�e���T��xB"�I��J�f4~p������b���M���c�Q����-Z�� �s����a�n��&SI-�nG���L3?��nH��#���1J��� I.�����	�����#��vb�}3
��SLK�����ٶە�A�f��)�?P�-Э� ��s��ƨ�'��5h}_�L��z�|pA_��k�����=X����T�F2p��^�I&s����:z�k)�o!��TDK���X����3�Yq�EC���
�.��3��ۣ}q���H�$Y���eL�����`�.�A����56���
 �\
�V�,�?D�ZuG֓;�E����D� ia<�c�v�A�I�5��c1��B�!��@���2d��%x+a��o%;h�jq����U�n���$zJ��r�[�w�)�Y�Bz��Kb*&��2t�tu(��8�D�®m�Jh� ��4�aSěg/Q� ��&i��q$�0�Fˆ�
2��Oƻe	
���]�9��g���Bc0P��v	�Źگ	
f�+l��"���ˊ����g@�������Ea�����Io_6A�^q���������c�9�.�H�=��O/��UB��Gb&�eH�9�$r^�F)�tz]���M���8�1��~���b��JX��et[��g��yί&ޡ�3�?�>�2\/��C���ۣ��� # ���?97g�˃��㒶g�I=��r9�ҿ�ß�} �K��Z�$�kM�� �������3�v�o��t�S�����4`-�B�l׃K��j�*��^X{��ߘ]�H^'IFG�~,\���(UރȜ#{NB�0!z��$ab��Q�j���� �?KT�zh���#���܄'����K�JI����O%GK�]��i1���ǁa o{J�u������\�����bܻ=@+q�N�Ly�<Wc���V��i"� �E���2��<��m�$�b���L�r&H�ì�nS�����b�ߍ<��{u��r�;�d��(��]qɒ�1�+�9J���1�V3�|�4��]�d��א,�iRO�����ڷ㭚U�~���/�5�����w�n��{�@�Mϣ�Y�s���Z���D:�yC� �P��g΀Z��QEV*�{����L+W<��Yc�ǽR�K\����odp9����nb>�=��K��Y
���=�R����7���CD�:5!�-�U�����~K��[�M2�v%��s��T�Ѡ���%��^���q���z�"Y	������d�4Â^i�PR�S<k۩d�xU�0���(/#��ᥧC2V9\�LA�U*���E������ۍ	�dm�]�>� ��,����67eTX8��^�-�� bXUXRY�͹ۦn*�"O�l[\�gR�;:��K��1B�����>j|����4����۳1�x@'w���D��_]"�P���ҡ^S��Ȣ��#� %�����u��3X���\ǲ�4���=���w����B�"�Ur�����e��jnv=_f��	�����Ǝ��_%����9��؎�tb㯖^�����&���/��Pr���$��0�X���t�}�>�sl��J��ᙦz,�g^��"�z4�`��3Dt>�.�d�$qFK�o�V�����D��E�.�>�O鮇[�gH;��4r���-�mޯ�{�uyg�7������ES�=>�Ӏ5�0/|��(�*)-C�EC�;U3�޵���-飍�񜐛���.��-P�!���Ju���gq�։p��[Ȫ�t��P{Rv��W�x�,߮&�(��ZR�U��|[/n�%NY1����r�0� _��՜���G�<.U˓~myfi�^�� �s�b^z�L ��v�ڧj{8Q܉I��q��pf�cf&�U�d@V��r�k8��j)�[pA��op�� ����23�y����_�v卸5�<=,XĨ?c{����K�C��)��Ug���~�^������t�)�o��&�;�JV����^���j�0^�9Ȋ�e�K������8���A��¢8����T86F!�ݡsĐ�&tX�O�d́@!���ur�!�I��U&���q�\�Uч�T�G�5)�ϋ�-���X����6)aQ/%�u*wP-MB�	O���T/S\rY������<�W��v/r��b�>�.��P%�&J��5C�s�t�Sh�W9��d�>AJ�I���(k��������+)FB�GGW:X�b�o���s�nKx���� AdWᢆ��H"oZ�t�.�zPy�o��|wnex���zAe��1+Н�������zk����N�PI`�0�k���h�P}!H�쮃v��`���E7��4g���@��fXBH��<�����tu�� j�!�%I��������U_�C��7EHc�1*y�1���g��9aB���Z�'��s�qR�� &?u��l}���\Ӥl�Q?E-'�<�*7����L`v�N)DD��ǎN��WƆ8D/��3����K/S���n��n�LrQ�N��_r�Y>��)1HS+۳��x��&�4Vj1���b�8��x�;�z{��$xv\���2٤x����a�7}�n1�i��.��O'+�>'}�+-�/���/�.���
�ӏ����S�7MҬ�DϷ*�o/����='Gv���/�M��Z$�o�v���+Ir����mZ�W�K=%G�G�05�l���/�`;瞩[<�K�(�4>Q��s�8��p�c���$U@D*E��/z���S��2Ⱀ/�^���V\�v���ZZ0Q�Kaz�f�$���� ��C&^��G�Df�ҽ�xg�Ŝ�\�F��=�>���7���vc��a��G��^aT���>!9į��N%�\��d�g-m������j`��2&_Sn����綡$���XI(p�Y+�^���04]?#�E�NZ/PP�[Fv��ّ�n��^��q<}����P3�F��p��P��0���Z�ʣ,�vs�ў���;�JIȿ�c��>D����^^Q���M�z���ʥ��G��������(�f/ xи�F���n(l�C�ڇZi��m�Y�U�H_~�3��Vb"B�t2��sý��]� Yq���z�|�ȗ]�y���(��b���x3��1�W�XD�T���B����3	����'h;�*���'�灲-y��泩S3��B'VH (��b5F�#������;���tU�fNb��-w3I��U��+��Q&�P(7\/�a
�*AÉ���6[�|քq��"̃d��x�[Q�v�)k�c1�"v�����-4�b�����&Gl��H�������^����b�!5xB��  K>=��/�������W�d8�����b�X�<9�R&�*��4��ʩ�:8ԇ$ �
�&�� �������=��a�"l�	���Iu��� X���(3CI%XzlQ'�GT:��m��Q�wܠ
���c�r�>K�(��G=�HWk ��@΋ ���[}>��n�g�Qy�ˌ.0:��G��A�K�o�z��[�QG-
^w��r���N�P1;9=�E�<��S���_�.�Pd��)Ev{���ʍ}�eb$(��6��3���N�lM��?���B#�q@��{#���5��4�&���]|�Yv��C�W<�L���
�/ät�+D}`���Ȋ!C�Y87'�.��S�� R��7�#��/U4��i����Ҍ���h�o����oh�Ո.~�HEY���s@�K9���1��t��4̕Γl/G��X�LL��X�^x��e��1��FE��E����U	4���?��M�������<^��e�&u�49p�xU���@��.�dN.aQ�Fр�?1�FDRiÃ,*������A��C�6�F�]�\����������_b�<�wh�I$A�����x��<�K�	���C�\=�������'[��G�0Tl���Z�y͉�>M�0�S�V֑~�Љo&�l.B�*��zF6���W���Ɗ���EbP ��٦��@����ұ�_�����Y�J�$�s��L	�+�<��f��|V�i[H��[��*���įEkp���^f�������ۤӛ����&_�f�V��({�J�T�����%����J�*C����x�|��vS?�Op��+�B���sOS΋�Ǐ�j��'=y�"h?�ݬR��-5���G���x:�D�%U�����(P]A2��1���R�qkh��s��V"�;�e�6kv5�����Jz��%E}�~�J7��-5�Ѐ�d���q�!(���_�?L�Lڹ���6P>�l_Q<|N�U��ݼse��9F{�<�n����*~
čc�=����E��x�*�������p�ܻ��=��v�Q�	�x�3��7R��a,�X#)��/�B���L/YV�2O�s8�%�՚?,�\?p��XJ��"�X�laH6F�좪�(���Ӿ@��M�j,g����<��'�/�#u��H>z\�T���qk'V�|�Ei�ˊ6�/��=��2Σ�}b͇É�Y���Bޑ�5�V���ml vo��H��N8]� W<��]�ԱxZCˌX0S�4]Z%��H��,��s��哴���kP�¶�U����jbG���L~Cvz>$�Գw���e��H����6�,������ #�w	�AfU�wXT���;�u�Qb�6��2Z�6��*� 7�g�{�~��oo��B����<��D������F��n|(�p4��:���8<S��O�u���o��Jv�$v�����<����v�E��W<�Qi����T[D�YS�%�`O@��鹓� -d�_��C|���� f`���
�uP��.��O�m�g~����� X��1�ge��xsFt}��" �����\�Ä_�g`$F�=��/!�E�.α�[@%!���k��t�i�ې a/g+KN�s5�k�q�ǂ_3oP�w����$�V�r�y�,ZNv{T��)�P�ӌ�@��Nh nǥq�`�^�D�F� 3�}t�1��qq�D��ȵR&��!=���4��l�,��#�E��=�zG�7E<�� ��
%�ۏ�w�H���2��5���ae�y�}�X��LI�MR���/��6�|u�k{L[v5�H��O/��!$yr���V�ɴ�	��yS�*� m��	yn���MFVi'1h K)k_N