��/  v�d=<� /�����]�<���9o�I���a�
@�ٯ��E���j���<�CN��Hr*��7?�%�����d^S$�0���<SG���0}�q�hS���.o�o�X{R�?9�x��ּ�@�����Y�v.'1t��>�1M=�\,�i�R5V[d�v<��m���X#�m�o*�����z5�22�8�G4�x�{[��IW��(X(_<A�&��աW���xίe�A��L���*�3�����	�qʖ4B����$�����׈3�
|�C�o��D(�H�A���e��tN��˴s[��	$]�'VӞݦ�k� :UטK��Ǟ�H� �a�C��|�� �P�Y�v��K��b��g�?��w� 1)��9Қ9��}I,�/{����OF#(�����\x�XCמ'�è+C��4L�6
�e6�"�}�y�!�e��)��ܨ0�E;��]Q�rqR9ڥß� �#�	\�7�B�b�H'�jbd�P�2 ����o66V�-�����q\��b��0��)ϟ�b��#᝸�Nf��-�d��'��1EB��z��AJV�@}"���'����z&~\�8��,T�ݴ�����X���}�G'���RϢT�'E`[��%�e�(�qXQ�6�B�,����]-�/�}�M5@G3��kv��qO�]�"B�Լ+�{���05��\��qc�K��{G	��*�ZqX� ˷�x'د-�e�iD������������5�V�ӌ*��_�(ݎ���~��v���HGV{#��v6R�
�e�hn��{]�,���FńmY\��'l2�ତ�,  !�Co�@��&#�BV�w��>����îf���OH�]��d��mk�a�T�0�I�s)��?D��ײd��lUyw�	犀M� �tE�Im��@KI!�d0/�٫\�j�Omm����S�bQ�G�p�: ��Eez����b
K������g^Ƕǚ���`(kM���º0��>]�t�5j�,H�G)+�K�Gۤ���ϵo�to���Z+fM���n���T#.�Z��ҵ��϶ws���ֺT�2����!�ځ:�V��'+�k�A�S�͂�O���YX.h��KX�ޢ|\6���Q}�}��^Δ5!�m����*��:Tɲ�#v��� �=T	K���M�я�#���Ju�/*k��o��jᕠ���F?R��q������8�)�BB@��Ȥ��Z�1��F������{K��#d��`�m��&yL�3�����Q��r۸v�����.6'���K���u�V�hr�N���7��K��s�- �&�9���Д6qbnY�?�$ӕ���-'`��a�e��p����{�{Ҁ︯��'�Ph<mP�$�mT,�ְ�Rq��N�9^J6M�H&ʕ�����:
�,~r����SvV����Ep��8.�2�# ��L����/�|��&��(-�䣻�Ѩ	�?5¦ [�9�'{q� z��v.�f7�խ)9��J�C�y�Q�t���F.��b�h�z�����ZS��4s�ޖ���>2���*.�ٿ�Mt�$�u�魦�%�7�2nw���s���(�<Cv���� ���:M�0(�֪+M�=�<���Uv(�%eB+9�s!��pI��=��)�frSֿ��-
��FD�X���`I�w��C��k+���qC���zUv��v,�GV���i0V��r�*s�Pګά���G�e��م �f(��"g'�8�E���i�V79����E�]�Ͷ_R����~�K5��r;{i�����\��d�k���e�ӋK��2��>v2PVѾؐ|~���Q=����sC�TjZ���2�}�U���Xhy�O*i��ԩ�GK��l:�s�s���z�p��	g�:�͛������:̟�C���5��ޮ��p/j�����k��4��2�%ZX�u�X\�2&����-�fdd3�m�<�$."@74�� ��ό�gП�!jg��S��Ԋ�X��Y4��}����2
f�[�6�6��g?�D߅ȴ?;5��*Vi�&���FF��Ӝ�\�E��vrlI��H���ONmX�ɬ�:l��f8ģ ����
J?^�������tI�Z�3����b�n�}��{�X<�ɔc�6��v���|\��W�tv}-a�.�3���HAv_��Y�v����Q��G��9W�ݺt���d��{k�b/v>k҇	Wt	�������Э���,���r{#-�� ���H����b�ua�1��#�	�R;h��g�F���Y���QW%������&�}*X�S,�_?��9�;���*`aGZt�۟%�15pbzH�|���Α�&W�ΛU������$���]�f��R��*9�pI��\�M��zy��o{Jię>c(7h�s_�o<=g5��Y+jV�nu�D�+������.�-�y�0C7�1K)gs���4;��揠 ӜtO��j9~��A�
�?�()��D���Q�Ө������43��nWo`Uii����:o��������r8fp�f�����&=����4aR�9�����{�v�1i�E���Gx/ҿݥQGyCԒAH�ke�q� Ũ7+\t=? ��F���3� ���.2��"��|�0����nM��9=p�
��+�S���J�'؎z��{E��t9�R�b r:5�$�����ņtq�c:	 N����4 B�|���1��)��`w�n�g�+�L3ʬO����ᙟ���?�����t�\%j���!؋����y���/b"{�lg[�!{d�A�$�뿕c���򛬸��@t�͗��a�v,���q´�J�,	M�tw|L��+���	�q'�����'d���D����"K�w�nc��܏[�fX,��}��L�ùn�m	M���bt���$�]��[�
b/���1ݺ�
��
��⣝�mj�Do_�B�u��G���I�E

(�qg�J��
��U��ZJ�H^od�Վ[�2D�/G�"1�$['��mujPڒ���|��G�O%��?�������i�,#����<�)˅唩�v��qS(SP4�㌡�An߅Β�x��"̓���=���1�l?	���:�Kv8�"��o�V��[G�P�ıe ��-� �ƴ��+���nKeʣ)�-z�5<<� �~+�-�H�=�����ƀ�,�,�L��ћ����q�
��?�"�j[;�y6��t������p�^6Y2�����ʯ���� �C� )�Yf/��re�C; ���{y���w����~d�uʹ���J�-	A={�
�S�L�1.����d�������\���O�A[ ��U*�|�6���b�ѧ��e��yiH�?0��[X�px'7cg���ڊK靪J�e��>Y�NP�ٮ�FaOh������͌b��c�FUӘ��9�B�TZ�I|��J�&H�=�E{�����7 +�@gs)�o�07�a�t�A�s�q_/����*��þ3l9(}i6:��(��y�ڜj��M�� [��^n�>�E-�گ�TH~���;��}I����ֱ.����X����	�4E�A�D1E͔$�V��;� ŴPLA�]>���Y��3
j����Ym@����X�鈞��kQ�����ͽট�av0�S�>��;������rPZю�Wճ`��|oRk)@6V}������%��0��I�l,���{� 	�.c�D%��j'"ڏC�f�7���h�6JTK�z*�J�M�?�S���z�[�tbY�ȉV�@���N�x���C�����Pr(^�j%�d������ψ�l�a*��L���ښ܆���.߹�n�@��$A��я�F
�F�3��Q�Ю�n�{���(�*u�_.�����yT#{�k�l-qX��_Zw����a?�S=$�4"����8�h4HS���i�Q�k�_i��R�̍�_�7n��v�K1�k��Z[/�T�&;�S�/����R����i�{�4�5H� �� |a)�u��.`=���� �b���e�]Gj�����}eN��GJ���D;���ʸG���ʱ\��]��e�$8�:�֖K��\��~��Rg�A���c�q��Ǒ�Q󖚈���j�4X=���:���c���N.�yC�Az��C~��,H��*�U�4�*�� �6��V�}p��M�b�s�)��2.���=Q�����"����2_Б�)�hK)2W����Z7��TM���9Q�%Xͪ�Œj)�=��@�{��+�<�s���GU��"7���s�[��'4�r3�{AXH�� `��G�H�ݭ��!�(���\���b��2t�`n�	�����L�Y����/l�Px��'{�!yM~s�t��^�2u?�6���ž�wO�B=�֮a���Fv��l�ז�X��J{�f� ��®M���0�Cձ�$���L�'c�����Ɲ�oHUa����" �&��n��:f!���NQ3��_ŷ�������qǸ�r�b&��>�)�4���*�}+k����!>���a��E]�~�hW�x7��[�����Q0 2I	�̭���fa�Ȉ5�`#(��͂OZn��U.`�����2�|<�����ar�YI�W_��r�0ȉl.���!��%~K��E	p�%-�jN����O��{|�?��;J��m��������ӇAD��3�y ��#�ޯjd����	�b\"K�`�w�%��+��d���`�_��(:�܊`m���ޢ��5�BRQ�k���v���A�"��dZ��3����V��@�(��o��M�Ai���ŵ�\<ē��S�(�/\���7�	ggBR����Ft�����2�\���*���B�2E;GE����ª���1���O�bw'�!u[>/��9+����D�伅i���QHs ���<�C�������7�,q�c��}�_�X��
�%i�Eu|�,�{bK܄�S+f(�&��s�X��/�� Ұ�����[m���Iݘs:Y�b�_<��`*U�lRI�s�g� �_����/���	��c��x���.�8P)�?��`��б]�G)F�z��%0O���C�-9TD::{㉅�"f��􂭲xI�r�'T1]�~1��h�z��x瑔h#/�2�x0�3e�t����.Q~�ދqK���]F;�P�V�s����0�`R��������q�-(U�@R��d�]�����	�2��B���o=�]7gW|V��v@,�N^,�i|�vя��iտ�$�wU5Ds�Z��z�n���d����S?��W���Hn���ٷ���Nx]Z��L](���bJ!�+r�ӕm���U�ؐF]ːvF�g!�	���̤w�o�_{v�y�OavlzІta l�<;T�A�?���0��m���������K��zse�����0��u�_CS����`���WU��Zc_Эtk�?�w�1�E�4LA��vA��G_��3琹��B�!�n'�)B���Ta�&c�p��1����j����V�`��,��y09�"�C"��҃#2�n*��5@l`�ȷ�E��Z���L�"����e�����n��vo��z�I�$����Tr<y����"�9�����flIA��d�Z%��z{#����0ש�jI��s���т�˲9�{2�$��w��b�P���Z�Z0t��9t}nY���[f]�c���l[eG-��% /�����Ti��yZI��t+I������Dxu�9�H��kj�6~pn���ʋH�R����@��P����ʩ���D�� ��F������Z��'����zE�J����Nr��ݜ��]
,��"���	�뢼��z̗�2��<�����a(l2��0�v��N2� q	�Mv�ۑ���S�jhKj����6T*y�X�Y231VXp��lk$�`�|v9�IË�D�xo!N�m�fx�L��wUҟ��?�s] M��1[���;�핰� EF��3�U��e��|)�^x�g9�q��(�v=u��!0~��q�� �5P���.X�oX�6|tG��Х�������1����~odzc�@� #���/E��%�w�s[K
�
�Q���l�i�Ő��@g�$��ރ�ねH���F~ɽ'~�gڵ�s_���<��=�������G�JymW��op]ۃU~9e�-��f!&D2�ӖBm����p����x�z�����Ӝ��R�7��"��xr�͈<�IF
v���D��XZt��_���	n{ۡ{�q��MNx�i�ζ��e����B��9�{ڏPK��L�S{�_����*�e�U���	/�wMx���o��=��x��KI:�Ϭ�ž~�l�u���l`�����r��	L��OY�Cݿ�Me�$����Xs�<n�J��>�](o��KgqhZ&��܀�~2�|��ZÎ��A���/ �c���:F&<E<2�Q�8dU���儴SL\���^/�Bi�NX�W 9g���KoƳ�z�I�Ge'�Y]���ޛ9/}���g��Q2������V��p�}���׹$��S�Â�b�d,��U���4&�c-xrچ�q��yB��c�U�&.��lhn�Ψz �Sɀ�;P:�Y��U|�w�2��Քl8��;vCoB$�)���1��0����
�u�l���.�sʲ�ҟ�׾�sQ���3"G�����o$=�w����ޛU.�R�@�݃p��#�]ّF/p4�T rF�p^*����:O��<��CG�έ�&�A{U]��w{8��ޛ�_BR�)�X>.r}v*xu�����n�u�6<�����MlC������� Pf��H�V� h���$c��|OF~�c,�c��VDRz�(���*�Wp��%�z�iv�NQH��\(�n;��}GL�O�%����]�9�{���-Z���)����?3��|������ĺ��*���6+=¼�/��i���LI�y��@��������*+�2�����b��"�z��_ax��~�,P�>�{���"UtZ�$Y#]��
�ƾ��X;��M[�N�퇼5c01�$kx�1��dSpϠ�7X/�-hf����x[O��>�@��x�ܐ̸��ҡ�ˁ�2u|���zÁ�����Z8:����W�5�A���� 8&�6cm�q���m"�x����><FBQ^BQ�D��K$�$n�0�ؠu>ǵK�)�����ba����f@R��������n/l<�ɁiΓ��/d!1b֤��4
�1zϭ�pvC����L��#.��P�m�tJ���<Dc�òw+�T��1���Sǧ:e�8@U������UlCHy^;�'˯~��9{[�( ��8���m�7���$6zw˻�nq�7>R���
�2P�aLA�XĊ�a@�m���ׇ�K��5�TA�f�&�#<$r��I	�C��W�\��#��#G ��� �x�{bET]rl�aٸ�0�=xKB�Z;\#J��8�&J�M�s�{�Or)�Xx ���������8�a�L�_���;�1�A�� ��Q6�����5[�qQ�G��3���%��#5��� I�Ǜx^��hǬd��p�T�hZ�]�7\]CJ�&9�%��X,F���'U|=��;�;�=j<���^��f�8�X4�D�?��)"7�^��[��;M�wyˬ��DZw�dܯLJ{k3���+���$/�Q�7�v.����؄�`�n Q04�^��L�U�RM�P�~��C�Ģ��)��&-�k$J8e��_?��x,��E������$9�4>iD+�|wj0�ТOa�����1�^C	Kq�����t%���������59�u��mטMH�E�3�W�_���m҉6�䥁V\dl�4R�1�|E����	���R�k=T|�k].ȍ�dG�5�1�'�N�;;�}�+F��pP#�� ̪(�:�!_�ĮcG; q	Qd"��#5Ҩ235��t�xp�:o�=v�u�z-�D��$�^,�`N��i�+��cWfd��3�.��Sf��J�H�>%뀩�F[s]C�lu�0bP��+�*W�d��������ƻx����f��Ki0�%�2�<o�z��0�����M_��t�N���l��f.w�J�&��xd�St�q]q�������9�T���5���y��0X�/�D<]_	SC��Ч�D�0��^Q������u�K�W�,�&��X��G��HH��]��O��K��ߨ#�q�<���_[����@f���T�ꙗDX����-j���n"P��e���xuaw|f�⿁y��}7��trA,�̙C�7�ӫT������� Ŭ�̨�@$��xϔ�	�����r�6����c�d���7,�a��n[�d��䧤يKٳ�NE-e*C�W��qO�1���[�2�c8����w�d��Z%�$��$��j�����l�2�AN�b���yPF#����	�����h+���/��rD8����p��7H���c0��e����K����×c�s��b;yz�ؙY�ql<*94Y�fߍƑ(�����̋UQi>NӸ�H���$��[z�Tׯg��%$�>�x"1N�;�]'���;7��6~om�����ӄ'�er���a~A �[@u|��6M���U�hm�r��<���)8[p&�M���'!�[�a�Ȳ����x���A�e�2iw����v�ޖ7Hȫx>���	C��|����G3"m�J��cV>~��D�x �G�Q���<J�bȦ>�N(Dr����S���6IeC6픬b���qA�����"}���1�/�_��v쇶|��Nɺ��ox�u�F���p�����'���[�����c2)�7,������]��f�3���]�qU��A'�nL+p��e�?e���y��T��D:��	nX��D�ISƗ�L#��R"�=-��m�����c�L�{Q ���#���7��4�K�ʮ����lB�һ��Z���M��ӱ��.���l���ʋ{G!~v5��"e��@��WH�!�lpRL�*��qm��n%��f8�"���"��N���5�V��O��P�*�fA���#��QZ@Z�g)�=��ճ$��5���Q�"1v���}���~�/�x>8����! X�q���d&�kC^a Wח����=b�N#VU@t𙑓��=v{�e�K26�$Ր�Md��F\�a����������`��b��6�%/*/�RGo��&��}��.\BJ5���r	GO�l�� n:G�n���j,Lk?ۏ�\����r�=��9��E ,�n�D�HP�S��&�hp�q'��:���M���Nm��7��j�&z�0m��{����̨��;���:b�*�U�`��ZGK2�F��2FCR�-v���}7��GO1�t�=�iHt��<_IB��=mp�y�8Z�#\Q�#~3T���#����Ծ)f^�[�X@��p0��ulg��>*㝅���^^Ui���ƶSգKW�O �X�3����{R�H���Y��g9�����uOtN:ߌP|o7�z�B��Y��Z�_�,|9�������lH�)�lV*Ph�
4�8�������j�j���d�9ܑ�	�(Ɩ�,�p+\%���;����VV���\~e��Dr�+�5�c�B2~�����+L`�m�V�k']�Z�c��Ew��&��;K���|���<u��K���X���nf'�+�`iQ&]ylSf��53�zs������K��=�X�N�O�yJ3�U�9�?�	�b��)��M1� �W]�/^P}����4 n�z���;o�m' N��#�������p��@��Q�5[TjSa�l��.��J�����Y_��?�	?=����T���y��z&-��[,�z��fbL��,4U6����ߢ1����$�t���u� )@4�:Ֆ�=B1��e�{c(��1U_Md ���۽=j:��8y�"�-�H�Ɵ������j��p!��u�f�}R�R�&%&��(����}��1(���ĳ��'�h�0T�K���7Vn�8�gr���j���	��z�t�T�?ٻo�'�Q<9�y�B���Y�3h�
do��W�uM���ܨ�<�4���Y�=߿&���4�ޱ��Zy�.�.�Õ��Y�S��YDK�Xg����rq<��j��t���U@A���6���3�Pd(}4�<�و�T�:�~�lI���X"�yS��z�!ς:`��g��3�޲��Pe7���1*����ƃ��t�l��2E���ztG�Pq��k΋�D�	6��ˁ�tNN�V����!F�VQ/�^Q�
�`Y �0�9��y=1�Ƌ�)���}���Et�MjA�&e������e	I�dp�oX�ܑ�0~t��z���{��@hFZZ��U�ݠ�֬*ꐷ�_	;/���~VI�U�\^7��F�+VӬ=h�tVq��x��qUnqA���!q�m0�l��4kۯ��a&�� ��(��K��%�S��ޫ�@ݧ�d����^�V7�4]4�����	����㢴=A���m�c=�w���qH�H����_\\[�U׹�T ��ncbĚ��S"�J�\(眘�p�TҠ	\�ѓj4�H�c�����l]��!�&��oҢ��at�d��?,}R2��Xȑ6�}�%+U���p��z0
��;4�Ῠx��|�B6[�԰d����2J��e@�#q׫�/�ܸL�����q���{���3֎�P����O�l��i?ro��K5�	���p,:XJ5H4�J:�>��D~:�V����P<���9[L�^t�z�t�i��i��:�I)	�_��v�I�6�}aP��"�hE���]�k����z6}�OR��}��h���t�����p��ٮ	��[*{r�4�i)&�@ɻ�p!;45P�9�����v�]�~��Ah�FL�=Mz�\�9XPw�W�[6#ja?�']�H��z����F�,^�0�>θ���@�b����X}C-��A>��,/���s�����4"V��e<����n��ъ=D����a��e�G�E)ו�HG��j{Q�Lk�+)�֣�U#5�AH`Г؟�JQZ�i�t4�;�Qt}��mr������EH��/y��N'k�E7YD�z��Q��崓�?-�*�:�vf��-&���� � A� �ܽe����F�eANf���V_l,)�9>������N=���K���/xڤ�1����	�dTu�����!�R<@�f=�
�6��c3�6ŕ�%S������1�� �Ft�\�I4�L�K�yM5�1���I�l�I~!:ms�Ch_�T��'U����<��l=>d�x��ϧ
3���}���Pz{vY�(޽�"+![bMeq�ϫ�t9:��we���t���c������#ք]�oX6
���+/�o���XE�x�w���J�s#"�O=���5&�"�3���I-h�f�h��ZG{��y�u����}2y�,������y�n���!R^e�; �پN��9��D#��|x�+p�'��7R  ˓s���25�	�5u�kky��1����^o�W�T�>�L��:T�����`��m�j�6�����S�O� ��jJ�v��Q��;�F��;�O�K[���7�L�� ��=�.˧��'Q�gx��������=�r��$0}��vN5#�$���RNkb�K��3-*+��0͍�T^��7����=g/ߪ�؊/����-�������!��#n�J�ʨ|o��AI9����e�������I-;��P�Y�������K��C��):�D&����3�p�Ů/	Y��G�)��GWN�aA�S��<�*�3����N����Q�
.,yѽ�=�T�O*�$ק���Jv��`��W1������S���d�>�'����0WDn���3knK��@�:f�5��j��i�^�3C<iB������Yr镒�B��PQ�BGu z3|x*��yE�
�X�/��vO�]��f{I����Ob������eƧӘ�뾌��5�v[��U��E��A)e�}�ҚUC�~c���YW#�qjr�a�C�qQt!�q���� �ȩ�q��4�S���,��Ji�$�������\(l���T�A%ķ{��l��J�{���_��B��rE7'�0��
����F#v
��k-W��R+�$�U�ުcд=����c�[B:Z>!�H���i`ʄ7�Z�6+��n���a�h����h ���"&��w�¢��KR�`��N\�N�-�,3o,R*B5=���眹�}i�{�%�8��	�:u�.\�"�:a��v?~M��z����II�qϩ5Q2����mdl��.C?z�T;��gӍ�Na�������j�\�BF��o9|E�"q�1&11`��O'ILU�X�������S��IP�X���H����|��^��������C�Q֦M��OG�Y�(�������وv�K6���ʁfK�Ή�7/��BqzG�:����e��xOmW@��?���q<�84* 1�Lz�p��]ӽj-F���íFF*�,�L$7�dx�/�u��!�8ÿj���V&�o����!����$��!cLB_ K�ⶴ3�S�ə�|��X4���.a�m#�$� O�r�E?�8LqyXIlw����r7�[��ɮj��cr~�3�^058\�!��N����0��'�r �.zr��� �_��5��ʽ&;���T�S�o�j/Aq��I/����y?����D��3�&
�T��{�H��D�����UO���84��(40�	���E��QϬ ����#M����d�1��~)M�P��R�^W��k/��j�^� ���dM��
A����=Wi�ȡ�6gt\
S̟a�����S?�܌^x@z���,��3�.���2��т.hEiS�����v��r/֐y�w9/�H��;B������u�=*M�
��>N�yo[5:Ґ��WRH����)V�J�����Mbb��@	/�H������{�O�O��u9���Y:j�{����9٦@
!���XleN������{�Nq�%\���˫����-<�n>���3\��-���:�b� ��x�?�$�
��{��[+�!��#m�0ޢ�����9�"2a���+׃/�I?��h �� ��ȷy�ߥB�����&�[jYVVR�,Y����7������Z1[�u�T=$m�݃���IJ�sF�)����W��	�cX�q�B��s�^�G��ڲXN�~���eq%(#��d����QA�rT�@����'s˹���0���br0N�Y�L
w,I)�np��U�3�dm?���	ƫ pG�P�i����W��}�#�~W�L������`������Х���&�.J�A��*��]�i�UBV�+� �2���3!�5�����Σ�.�AX�J:�K ���"�#Q�-7|ͅ�f�r�q.�T	= Ā�`�?��~�T%ڭ�?5|*�vȂ�t�����ؘAZ��4��e�9�S��ڽҨ�n�a�C}�fXW��iw�$#T:vCʪ��,}�|�����d.>`	P�V�Z߇꣇Z����T��ʨ��K�����ah�%iF�w'˯<,6��N��Ta�,������9c*Q��K����ߧ���la��.ڢ!���Aq�w���v}�ŏF�㙁nO�l��JWjv�bh�6�,i3�Ba�붆�u8 ��:�7k;'.]-Ek�yN0�=�dܟ�x�o�zcP��C`�������sˁ�.��]��7����H�r���w����j�d��Y�r��:z*^5���T�n>8�E��[�[ �xBa����ت�5%@n�x�s��v��,M-��ea� �l�q�N �k^d�4�lL`�*hG�����Q��-=4:Z��|�-��]�7���(�Z^���g������C)�b}*}�U4��������Z�v�|~���Q:�_�����YޛZ�`���'�yF�)D�?_���ɨq����AM�Y�l���Ng���Z��.�{/Jw����}�%~8(�r�|����싧\6�#����Կ�l �s���E���J����N�2�cq�5D�KO��'3��x�z�C���F���b��V������AO��м1e��'��Ru\P>W#�|ܥ�)
�C�Ü0�a����}Nz�
�)���L(!�
 ��\���|�5!�6���/T��1�NZd�~r�8q����a�#ٹ�cx��f긥��+r�@DTh�h7���Wv%�N�gNB	ar���۳�"
�3_<�'6	t�i�cgnGh�j���0����}+5[�69�Y�	kM��<��g2�LZt�Y4�;Q1ё�n3�����
(���sX���.eu#��j�h�#$TF��kZ�'����OZΚ�=�s�GD��q�qv=�O��R���9NIsW���-��]Փ��L��>�~8m�K_TF֧W����ʙS���
��~���5z�����/����e)GMW���`+S8��Բ`0f��sqtI���e���u�:�\��[�YMb�\9�kcbV,�`�W����㋮_���(����aAΌ�l0��vG1"l��ax"���{���}�K#~r�@j�'0�_�aQ�~��P)LM�_[T)����=W�t�d������p{�3�i���c6���'\]�f����-2�Í^h���)�-�PKIi��K<����A�Ĵ���������"*������8�]U���a�N�1�}a���i��P=Xt�!]B��)d��?C� t�;3R�<�SԚ!��Na��/��ԅ[�pf�.{;�V9��K<L�Lى�K8x��hu�޻��kr�F��ʥ���L�"!T��K���t
)�Ľ:��D>t��d�-����\�1�֎���I�W�1�X���c�Å����Q�a��.Z	M\�\ǆ�Q�5�Ϧ_�'��> �i�w�:���=�n]��o��.�T����vbXw�r/p�n�=B@i�]/``��Qe��=�����gך-[$�x��ƕ ���Nu��q8����݇�W$��V*���WSM�S!/�g��;A��dP-�Wq�OBP��VeG;�V��P�j�鏿XL_�M-��Pt|p��P0�P7ʦ0W4�7�2�j$
��ߴ����& ʽI]6<bv#��3��'}�ܪs,���4��H��o'�U��_�N�;��6E*�㵙�6�K�&S��U���%����;R�.n�	�sV܃-�dJ�9v*8~�#���3.]�6�Í|�z��uA��ӧ�3��2Y)�֧��d%�� LG�]��1a�4�`���,��ǐ�yX;������x�&� ��v��7k��xX��d�l6ٔ�6�Ï͇[�������]{�*tpz��M~Du�����%ΐ5�=Q��W^��O�E;���4���{]���qO{�~�Ԋ��=��
F��J�<؜��	ڝ���'MRL�w"���}�i�Û{4�-�0�(��1��[�E��	5�%�����i7�H-<��p�
��l��5#�������m����]�6�m4����]���@���%��cI�4�=�0�Y0�x �ȹ��Е�U��X�Sz�R���+ڂ�E�G�6h�=w/���2X����_�)cn잶I�n�%�rH���px���e0a�R�x�H�%#��R��8�%�܄sR�p��/{�vl2�H/�	��E��Q��d��|b֖:���wk��\AU�Hb<����Y�ϴ_���E��O05'�X��ȰY��u��EUI��]=r��a������c�b�	�G���1���Bt�s�H)[!����mq���p滍B��t��	g:�$�i��Λ����Ŝ�L�}�qa�����>(R��t7}ru���W:8�����LT�FҴz���Yzeb���~�]�S{������}��MvŲ��o������`��w�iն+Č���J�固���`o���"�e}�N^ �W�o��g��)����^ADӠ"��k5����U�X�5��/u
q$+��m��p=��s>�X��(�)E�J*tv�Z*�K��[��!�V�C'��c��³�G�r���@�3��Y�<��ETDu�нP���8q�:3�������5�<q�^NOy�d��8�W���nZ
a�Y�.E�+'ql7ָ�d ��u ����d�v�~􆅗�U���-MR�oS�w�o�'X����Ց�x^K=ϟ)�Қ��w�nw�/� a�K@X�6rM^6#Ύ�$�;J6� ̆f��F���J�5�}��Q�$�f��v���{wϟ����ݡ �s��;P����z��KbcJr����W!����� z���	z��~_7ȅ��1�e�w�J�#@7e�>
��
�{�j�n�)X`�C��f�9��k���$�Z�$�����|�Y�������f�N�B�\F���D$�������_���ن�~=����NCu�s`h����he�:�Ņ�]��Jܞ���p	Z�El̃��Y���NGZxH����V�p����j��9�wJq������jw����qAh׳bѿ�WOil�2Etc̽����;�(�:0s�^���6ø�ˇ��U�E��V��A��ηQ���YG�p/n��c�b���� z�T]g�մ!7|�Y�c�	@�zd	���ඖ�^�ѕ��G@]�Υ�]�8���e�J����@��d���]��%;��������'��`�s�B鑖�C���V	_hILC�+�%��5	ۙ0W�NW�7�iFt��EO�^O��IĨ��#n�2�� �, �'^�*�)4��r��*�B��m�85oْ��n������G�z�9��2�\5�H|.�g��,����!(���NK�Z��BVBp�����$<�X櫱Q���ĭ�}f���Kې��4����e�z"��h�c3"j��)�m� ��nz���\	�����_�i�g4��6ҽ;ۓ��K��K4��F�o[���U$�*�����l``(>�\T%$a�Ru���F�T�m\�d(~/�A��TG�du¨�=w���bP�S[m���$xPwwM�pW;t��(鼠��9���K����ڦt�Q�?*OxȚj:��]7F�R�+�4�󱷍TIe�s2�T�B��S��L��'��{� P��̸�YT���0���*��"<���b )�d@X����p�N�OS��*�2��<2�]�Ȅ��rxc
&|NC!�;H��Z�x���0�1tpF����ޙ��B;��&4(ӿ|��ZA����v6qRV%�}��TH���K܂eQ̓�*�S���p��]>g�#�P���G_���`���YQ�?h+�Q�mXo�:�j^��տ���	�8_��'V�\!C�2�r=Bb�l��c{=v+��Dm:���q��/vS���ώ�����[\>\(�tg��;�,����K^&U�������˖d��Im�V<���) ��hl'Ut�`�i���@�h��[�\�� QPo�z�,�C|;g��fP��ɋ��\JC�cu���X���c�6�{��Oj��Yp�Gr�/�ڴ�)ˬ�;2�{ЂN=F����KD+vt�9�È�
R��0Ê�O�/���/r�O�+��#���쳸�wF���``|�� �əx	�Ee/�b�ꋀ�)N)�ʵ?�-;?(�׾����(���@���� �O�>6�[�e��&�i=��U���r�S�`Ȑ�Ǔ���|��|Հ��HR.!��ηr�<;��p��5¨�ʉ�{f�Em�C���پ\���P�iG!H��A5�ڼ��'�J�����@��=���$�!�G�Ƕ|��5ep����骹4
�!�9���F
�W1J�5�۰S��=%j�:�<��$[%��QV}Sqi�����w�-�v�(�/b���iu��L�	=�y�S{��i���e~�T��71��ZQ�BZ��D
����B��'��>��d�p��B����.��g��f����(�wP�#�Qr1���+wG �Zs2	Q.͟�Y\�;e�^˞I䖒�Ͼ��� �H���;e��/�Y��U�Ɓ\�ħ�l��ݕ\�ڼy��A2�`���R����Xb>�H�rp�5]/.�UdEk���vI[X��h@VL��#?�lq�S��^��s�����W�`��(-�p���Yd, H~�CH�1����y{4��W�%�</��-�_���[�^���7.=ž���#1Z�A��4�t1R�%�^�0�|@����Y2�4�N'&tZRj@���Y���Z�,�\j�#�%ț�&����F\���Zߚ�ZY�Wt@���e���4uF��7���=k3��	'^G��� ����{�Ũ��P�̘i�������,.�;�!o�zRpc �g����;��cg�Eq��a��0� �Z���*��l����!?��V�?o93Wڬݦ��=?2\W��'���|��[��i�$��p�0<8�t��?�W���p�/|
c�9,#{��Q}�|R�~c������׽���"�FM�������X%>Eow�w��"��ܸ�m��]�9�F�~?�F��C��9���h�].���cV���=�t�*mg��|? u5�|�v����r�߁~�[w"�@�$�[S>�S�ͤv�1l��2�Ѐ<�B�b�)Zx��z��˧*&����Fcx�[��l\}"�I�|]�ȣ���8%�Pt���j)�'?�3�Z%���FH~�Y�V��F̍J��QG��`���uS��U��&�B��� �񾉡�������"��[^��V�9���q�:�DM=����'�����y��_1�c��Yw�����+�X�*�%����w��8D���\:��XpTf��Bg
.A���6���鈄ctR}s�Úp K�שB	4I+��%rTmJa�7�q+�K��{mq-�cR��X��:}b���Gb�z�ϭ��BD٭���Rxz+1��i�p��LAqaA�����e����^��ù.�J�u�4�[���!H�����'R�*�8]3��x�K�go�M�������~xܸ����n_.ؚve՟�8���+�Դϰ�eu��k��/�r�����Vk�h��ԗ��"�]ZO~�������@���ԲT��]��َX+��.��dz	N���1�ƅ�vԪ	�7�+��*Q���j���;Y��K�1)A��� )��[i�aw�Z=b��9U��xw=9Q�̡��&�ܐ�!��p0�7�,�#�[�?�m�#2}��Σ��2�'�,�b��Q�?0�4O��l��ZcWـ�Q�A������+?���%t���2���_L	"��1��"g���f5��d�V�n1����g��W�L�W�2e�t�S�t����HǷ�;J̅����7	m�����ʹ��{���xe�)��eDA�p����?D��O�dxF��)���^*�U0˝��'�f��*��SyG�q${yǊ�gRKJ����Kd!kKMA3��+3~=͆�v�G��h{'���-�5w�Mz�!XI���6f�M�l��/�A2��kLR��g��넋6t��k�̌G����ۭ2'�E�IiޚOG.0Ջ�}U��zԌ��D f1k�N�>�.�~ⵃ�^$��8�C��������s��f[���t���ľ�q\��'U�� 4�|;U�фN�D7�"A·�I{z�Ζ������+x
��`K�5_j	d0��ܯ0��tm��qo���?�)qs��Ƀ��{��ܿ�Y�P5H���S�~�I'�	9"�"ǩzErr�q
�ђz���P�,�5sh��Hr�y[S���s3��6n��4�_��rA�A���F`2<y������[�W��#��a��>���2��q>�,� F�Ff��B".���-�B�r^\�q��(Q�r�E��&��M �6$�^#יb��1m��U,Ŵ�'�aj��h�+l�JN��ԨXɘ�?p�a"W��o�\xc.s��"7t��N�m+R�'��x����\�g돔��3�U��~2>;�����pi4���c��w����	!����n��ɱ>�.g����k�R��K���a#Р,c@��ݱ9����E+��Aӡ�x\BUY'�͐��)�d_/�0�85i�0����hn��{���a� �ʡi�b�`����H���
X�� ��wN��V.9QW�v�2&-?�>�"!8�»o���$8l�M"{����I�tS�,�	���ǝF���,>�A?��#e
��.^ ;_@� :��Q����u�|ko�=<i�`�T泼���ʌ;uSǹ ߙ�L��'�t�L<���]����������n̥��k�Lf��<Pt�ŝ9TE	u�$�8Q��<���,H�c ��-h;�i�SpD�f� Gs�о0I����Ʀ������l���6?x	�������7�6�6����[���n�����8k�V=�D�����B�҄����F:?�"\��C*4��P{Ɠ5Y2�
Ae�9EڬD�ik��(7�-�g㺣��O����N�K'�:��0+���$G3����ef�(�/�e_�M3သ�o��q�y��̜�CS�&��o��$܀Mg�3=Pa<�NT{�,x"㺈R
M"&f}PN`Yq�~���WƬ�M���r���B��>�oCA���t乚ʝ�TPX��"�t!��7zar�縹�K�XX�� %O2J�Â�^�]���(�7Ѷ�3U��+�l�yyCQ�*GU`/���F	mkNJO�a���X�:yt<4H�Rr<�`���u�W�poK~[=B}fJ$3`U��~�Ψ�5*�:4i�Ϩ�ߨi���F|���49�!�Y*8c����9�hrJS�Сi�3L��<̴�o 2���kN3&a���^���ڡL�}r�h��k��~��E	bhcV����+���W�8BV�����9hn��?累_)6n�U�FF��*��N�ӿ�yY�G�K��[�����K�.��p��աS�o���R>f�$�3�TT�@�Q��G���v^�=��]Dͩ��T8V��������aWF�W�CG�G���=jse0��ۿ��Q-]�������La�YЉ�ǰ����r��F3���J��Hu��F�J_����L��J��z�Q�Hj���&5��]�4jK�ڮ�^{`|�avJ�<�k��5$��3�
��CEn��G^��>�W0�X"�a�,�fZD~�!fk%�,�s�9V��ƭ�c�r>>,.�����;D�>	<J���to�uE�9s�[��Ů��r�?r��ݵ�������%����dZ �\̏E}G��R��}�x��������uL��+���81bq3G��4nNE��Sx:H�r�N!Z��@��}�j�!�Ov~2AJ`���v;&m�g�ރ�5�$�*h����ɚ�*-ql��<ꮰ�@8:���y�OF�V�ڂ�s>ac�N�x+T�r�窝!H{������l�φ��6�XÙ[>R����v��]$t�����-�V7qV}Y���ЋJ'9�b<�F����9��8�ʾ.S�-�>�����������LY�M�m���c�=�7�>'�gcvU�p��U/5���+�I��9t���y�����#ʾ~��k�<��jF����S��@�t��^���F�Z�&5H��-�2�z�Rݱb���8�;Rd�3`��P�I/9.!�d岑��)�O�ٔZ�fO<SbH���&3MJ�X}��l�}e�K�dm#��JiI�G�	��Y�AK����Z�;��۬N�P��YDp{N$�S��0��Q��7�e<�1�E[NM X"K���2o����GCT�Vq�`���~?G��C�'�K���)$~�y�.��|U����;�Z)�&�����i[�lUrx����R�&ݒ2��� |�Z�D��8JE��-��9�8Hf;RZ�@�Ɋ�CRc��ceH�`�r�^ۻ\�cͫ�Nm�To��
��'�+��k��#<�R/f��/�{�+,]l�}����D?���H
�o��~:Ȝ�l8��J�F����
�z��Fq��;CE��t�G`D�يD]+=y�w��-����ÌD��s~q�w��CRD˴���bc (E�q8���s���%��w��gV�P�[�<�R+qye��ɩ� �^�s�nv�sU@��Y$LE+�~u�F�J.�7d����#�d-�or�UQN��G�SpOKhg���nA?�Y-��'���^JK���c*�	WB����GM(�c״�<�T����̣��1��!�$Xg�ui�*�Y���FR�m8�v�_��aAXD�v�5\q<R�קI��D$�Ý�x��txoЍ����j�JO�^&vl��@b�d#�4��9���ߔ��neLW����ϩ䥓e�)+��4�������p�z����,Q}�
�.�h�/ޭ��U���8�=��s���To��8PC��y�h��i�w���^ݩ}���~�8M���Ns}� &�W�2����x��~���no���o�pRT?À����b���L)(�o���G-ħH���;�a�o��$���%i����j�0�$��6�V bC����Z�p�\N�-�Z��][��L��7���mP���Q�y��	�`�f����K12^���%:�e�^mq֟j�-�RݠʕQ��X��WD���6`qT��琮�o ���i}�0�^��,Kl|��4`�u,+W���]���]ׅ�H_ܲ����HET9��
��wy$��'(T�_K��T����DD����(�,�Rt+���E�ǃ��������7��s�Wr�J�X�cdF�ק�=Iox�ź	��p�7�/�뭳���5�h���<;��/2>�̕��0����`��6�v��\�����	�������zk�ǌSC`>�}�;�~�jT�q[���_�����=�� ��N!�9��1�d~5�D\J��`%D���~(�ˋya3�#?{i�aѥ/��9�����`A+VT���9Ӂ��Ԫ�:ށ��l�a*U�H!��+;����$z��\���J�^Drx�I�d�g�9�~V�/�GA�\�$��F�ŞI�@>e:h�������ٓ�X�ց��7���]į<�x�_�b��v��{@�
�f:��oϞ���uM�6g���=��0X�*�CQ;���\�|~�����ӛ	��Q�+��L�̇��온9���$�࡚q�o����y0�v����]��drzJ��2���qw$�vBK��@����a��Ȅ��������`N:��E��X��A����A�%�/����&2U\��s��n�0�jy��t�WeB�9t;M�E��plB)r�;3��s˄����� "6\�{P��P^8�-5��9�����V��a��	{K&�y�F�9G�=��>��Ȫ�Ɏ6��	Я�yC�H�ޠ�UTA~�h�?�x��Cmm؋^�V��s�?n��JӞ�	�.4=��#e]�0*�.�RP��-�Za�=6hv�S�û�D�sKB绑��϶��4s�~��-J�ǃ3gI3�֌s'���w���������N�O%ۧ�5F�.���$(&0�^2�nۂy�~���G�Ԇ:�{��@���-
)����~�/;�/c�"�kJ�q���M)�\�}�/���Pq
]~5E�S���<�@��*���p&Cz||b�{X�Nt�PW�ڴmR.�]���\�T���i��B��˯��\�B�@�%|e������}�+�Z�خc�aoo?r/J!T����AW����%�4�m�iY�0�$�1
���yg��C_:�Q��E�9�����f$�k������8
9k���!��������̃��fe,l��6�l�Y��T��{ls�dπ�:��#˖Sɯ�p�������O_z�yP���U1h��[l�b*f���<�����jG�3�4����p�j�0�Nթ�-��I�/��^�6���Z�b]��Dl"^]Pt;t��*Q���pRK���缯�ަ]����c�-U��EE T[��G����'��틎
:(O��{;P�U`x�x;Z�X>�P�ҷ�ޯ}���뚍pH��>a��@�Z(�h�y�
>|T2�S��uJG�N�J�]1�m�q�]�"Fq�9:�O�_TKuR�����)�3ܙ��I�������p��>����H./w'��9��F�v)�����a�:U�pB�	⮰Z?�v�7GmrK������ӡ��V��}�{�h�h�<�!RB�w1
��3\�b.D��~)Dw�5�v���JgHj��?��z����F<��͠������������O�.\�Z�����I4��J�Z��/fD٩����>1��A�SDhCE���:Y7K_&2��t���;�4��O�ҟS��8���.�D"^��y�տ�Y[=UF�i;��$�i�#�5 q��i�7p�0�f@&a�e�%�v�^$���y��n�$���t�y����f���<���G���Nm�<D� [��\��^��LHn
6�W����`$h�1Ӻ(EE�o��.HqO����H��re_�P	8���`��q~���k�]�w`Je�bL�P����]Y�q�9� A���id���y�E5t'���/ͭSgܔ�a���~�����	�V�z�
?�a����1�2��)��*?ѯ�4��Gr�5B�bC��Æػ����̅���u��'�ę��\�CmE�D�Y(I�E��Rq�x�d7d�t9�8��@b�U.�]۹�ل��$�Q�rk�_'���5աQ�B��������U_��������ŝ&P^{gm���8��/����\c�̖;���a���?YP6��c���2;�HWכ2�6�w�6a�=ӛ�fj��Xu6�go=k�)�y�b�� )7��8Q���?�m�etc�:ď�5v�6J�J���˓bz��B�l]ȷ��a��t��J{�cyiC��[�|>��E�~��/���\�IE�����c�7 {�q�u��S�5K6~�+�r_O�c̷Ւ������X�?���N٠��\G�}��/Pt�d�9�ą�$=B��>\+�l@��N�g�_�qM�����pf4ca]KAב{Tf9$���J���]'���T����"��#�A�c�[��t���Gy�C���Yb�ID�q�׮��E�@�i��ʗ�O�<���D��>�e�T��~����gi,~��.�(� �}w��pQ��?�aj7x�A����'�7�2 H):y*��JN�)�!Y�N�<P,x�����y�����UG���5��%puM������"����&<��B}L_Z��$ �`����7�r;��0~1�$��vZɖ���vڌ�4���wM��#�2�G{�+C`��2X��K
`p-J4ǭj8Ar�L�|ӟ���x���f�-�p�Z]���N���=�Fg�������W��X���wP�(s�ɯg��<�,�c
�p�ߕ^ڰ�֧��@R�o�����3e?#^�4M�t �������G��s��C�3�<	�������`�}�ĺ��_W��c|ܩ� l������a2_}�YY���c�w��Vki8RT�6
?}-T7��I�����^��'bnt�1g��R�T��<�b��Ψ�-������m�&���J̧>部;���!��Ƒ|��4��F�C��[��D�{�a�Y����$�v�i�9��B�Ps���q1�� p��eC����'G�w���[_�O���G�ȼI6�#��t����X��	�aZ[ͣ\�5���F'Q>9�� 'uv�W�i��!�s*a.=��c�>(�ߨu�ctۙ�)��͚�v����$"a�?���=б�U%����0��� ��O��,�w|��>fp�~~7�n~��3��PL*P���C�SC�M�A,,�lI�2+_�����b�<8�b�s���T��m�U�ݶ�J/s��С��?,}�5��>\�m�[���i�9�]�䪚F�U!�墁L8|��q����ݠ��A.�s�nT��>"vo�%��d{�sB���w����J�^�;��[��u�J򚳯|p�NL�Fi��0�[��@�7�+1�T0��'tЯ^�-O7���Ȃe�$���1u (��(����Kq�j�QȅdA�=���!��0E����'��t�:��>Ѕ����m�5&7���P�X��*'�Z�{����<\-�����}6��ĭ�y�ٔ�p��˵�:L����h>?9�$ȉ��$��d=�&ſ�R�6������a��c�l� �GPG$��.���ϢMv�K�ԅM�1��9e�$Fbri���m�b�]���%��$���QϷ�4&L�y.�_ZC��y|�����)��Oj�JJ'귽�F�fP��]"�JWA�W���{R�@z<lAY��{xW@t�c�� ���lޜ�7�_�fM���>nL~�茍����&K�e�c���Yd�-T�0�i��2��+�\�d��,Ac�S��S7\I���m7���N���>���9e��Z�+��'�j����3G$��M�Z�X��W8��R񏭁AQ�`)E޻k;5tUY6�R`��yD�u��Z���%�n5��jx�=tg>1nl����
�����=��{�Jy�T�)-���;ѕ��D%6�{KAR�E'���%P���2 � ��.���_ݕ3O����_�5�q�ו�-/k3��dt�Sy��W�iMw�}.pi�gy�,1�!���u�7�Mnɜba-��D��fVO��uV���ʇ70ǟkT������h��n�S�����h��e=:�Γ��>��-=S�s��[Ҥ!=$_���FT�u�����}Ȩv��eg������g�赝l��O�C�8$��f�gz�r��ǁ��z��p|�(?u�2��@"�t����K�J_,�:^��g�!0�Ã�_�(LM�%�-3������KmH��{=�z_q�\o!H�j<�p\W�ڸ7Nv��!$�8��󾙤n�-���5#�4?R�jFY��\�e]�b�C�^�2.Y��L�#2��/T�F�9���9�cLw
S������W$|��Hn���y����gA�4w}�.��PQZ&��ܯn�V؝j-l^+7���Kn�2��Y��lpa�l�_��jf _�7D��
;XԤ�e|��'�C�ߢ�w��`��ҫ�<� Gy��M #i9I������qqq47��"
�&8�fUILJl�6���h��X� �D�#B5Q,���(���M����@BY
�����ZW��7/!��JR�qʝp� f�����V"���K!`��E����t3@�8�eZ��)�f2ss�>?cy�ԃ�|䡼3�w<���T{�z���H�D���+{���݉ptM��2QO5���~����ݟC"��NI\:���m����Km Ϋ����`N�Ӧ��'C�u񮁏��\S�iS+�|�Ό�'9��(v�)]ua3����T�İ�u�'F�V�m�˚��p���ȼ$/�B�'c���t ��_&�Jfұ\���`|��
F�Ȉ�Ěm�sm�d;&���7��!
��s�{���YD�����豣���@$��c��w2)���XD���7�3����4���%��WDߠR?��vX���D�fUv�0�LX�^F�&v;�O��9�g�cq�*�W�Ǥ���hC�VO�vi�Ϫ�d_�ff^�b��0ׅ���κO��^l�:�Vx/V��FF¢la8��fu�і��i�^�
�J��2�'i̫�t�v��v��u��iNI/$c�7��i
=��u�hX����$����� �7S,z8�X��[�����b�
�����;�Ԃ�.1�3�QP_����p1@�sD�9��u�Q49=V�h����J���V�����)�s0��]tb4����p��1$�K%�(_<���>"��n=#�&n��������
��3A�pXP�N������k����5o5M����!��n���"����w*��M��7Z=vf�F���[C�,&J�mf$�Ay&^�t52(+������~r�ᗆ6��W��6FD�&��؉����G)B䖄{�b%��̅x�n�a��˪C5� 3��nUlB:gC��n�VB�X��t  -�X��Rw�^�x�^�̶-��4�	���o@͆.LR�s��[f����jy1�[u"�<�%\!s���]6Ʒ��N��s� �_.�&ᷦ�W����ڒ�LV=Aw��o�`x���v����E���!w	���7�&����(�.�ʜ�R)������e\��C��>H�����.B��.��{v�aW� �%B%�����s��٪/K�����%عm|= Y�0�����۫ę8��L!���Mu��N����$wgȌ�e��8�)��9L�"��*���3f ����(J��y��ZZ������~
E�s�?��D�&ȼd��[�t�sS�B.wA+Q����1���ݏm�͝�6Z�SZ�i��l��k�v�?0��ʱ�~+Z��-m6��$��'51�����,����#���ʇ6$��I���6�r�0�3�N7��ٖbG>g�zT��';4/���rX��{�2R}W�� 7e��	����#X�+���Z{�:_�l
7o	�+�\R��~�_rAM+>�U�[�aF��M�z����X�z�r�o�d�:�H�hr T��I����I�D�u�Y�[���i���<�jҘ�d%��K���<񧉋*�n�!��b<�J�����֠��I����I���Uk�m�8}� �����K�Z�q�Gk��y���
V	��Z�� �{�A�]�C�3��id����P�$6�/�$L��Ȍ(T��bZ1�%�{�� o���<��u��Ɛ�z�!k�D�߾j�{0��z]=u�r��c��"?��4�%�4zA�y |ؘ�N����as&6�:�/���d��R�^�W<P�Ŗ/�����#��QE���Val�ētƾ�#V-;���%\{�eE�_A�-�����ƚ��.����p	�~�.����SJf�m���k���`�H�>��%�#۰�U��uV���~��Yl[�q���xɧ��{�D���-��d����o��]��W��qI���r�Q�� 	S.�#h&+�U�3�-['�B��c������A�s<Q��G��"���:�����lÚq��.��j~3�H�hY���A��8
b�'��XJ}�`��Aj����"�޼K�R���Q���6��u�V�W4�#�N��o�_{��Q	��UTu��z&7=Ɵ�V,���E�� 3����=�V�rF^�����a�1���t+dF�N���V@��?P��`*G����x���e3Vŵ��?Y�I,K�9�"["�/��:��r�D �xm4{�供ǔ�m�h��@�����i�֧urk��T V�����g�����M	���4 �? �C���[ȕ�.�B���/�e��������)������z~��Ul}<����!a2��ۋEB҂���7�U=�6�D�H��C�PT~��J�u�v��}���)�m���N6�a��gp��yH�(�� _��1T:����Ƌ�k~Fv�p��;����hof��4@)��y�=W'�q���J(�7�R�������0s��9pbg<�0� n��ڋ<��G�P�)'o�Q�\5k���A� ^Z�^�BȾL�Q�M�T ���b��Ý���A���ا|�]�Fr1�)���O5g�����8S��p )f�8�e9�[�%?_����F�jW����:�/#�E_36_	�]�{Ә���=2�Y�Xs��(�*t�Vds������5��5�ۊ@=�U�"X֛Iۨ����?x[�q�+'=_h�`#�&%RfR�(�!)�b y.���/ڇ6:���N�5�pR	�������e����>w۴RF-��� ��K�oX�R�:�N%�1�0 j�u�ø9 ���S����O$cK@0<y #��.G�=��<�BRb������[���H�m�>�<��E�w��@��CJ>Ƽ{����T����!,+��H�N;!"����J4J�ߵ�7��X�;���y�}�m���m���	��X�����]�q"8�z��v�\�|;Ǉ~�Y��NW>԰��2�5^� �OҦ�L�4�u}=q(~-���B
NA���ΐ=6�S�	��|z��xr�*�����ٻ
����(�L���x�~�����նn0�kh�����r26ӈ'�5E�3�[�}�=sb'޴i��[�IOP�U�K6��Kn�K]�]��1<�x�J�����z���I��x���31B���� ��ѯ���LU���W�0�������?p�<n�D��������c�I� ;2�|��ZJ*�����o�A?� �.2���� ���?��!�&v�����Jc�`�����꒶��N,W1��Z<7�U��ń���'1���e@�-�#�ɠ��\�LS�W��W�V�9�$�s�O�ΰ��v���z��H�w,����*�V��Q�^�;�=v�P�7���k�_:%�*hҾ'���^c^w�k��p���Y�c�F1���s8��oQH�I�I%�e}�'���R��/K%��M��t{�)G���9������T̆�
�����S	�Z`�����d�.Q�z�0=ԪH��:�c+1�Z�B��|_{t��w����2�����(Q���!}�v��iۇ��bd1�����8�Vl]�2�G�gd�$�F$=kP
|�����O:�P��h@O�8g��"��Ю����4�r.�#��~�U\y3������?|Eץ\ �P�LBd�ɷ0ݑEڂ2�a�v�`�?��
%��4���gIv�k�k�x���u8��;�#&[�!z<��ZS�$H�k�ՍC���ߗ-�3�&F�����V����Y`��ї�� vG�o�8�f���k�A:�D�kʁ����0�:Xm�x�`,bm!��vZ�.�{d}T�h$�aӗU�lOV>r��8��ZV�'��T�.t��\J��z�sL�H���>j����ZM�=��@�T&1�
$\Aٶ6��P�^��`����+�De��:g �)��׭���;Y%����%���v��B�=��]5���
�}��?>�}й��Ή,3��]I܊f�e��Pb��x��@���ɉ�>�%������mxD��Z#�t��˂��G�,wS:�UZSW�^��W����A�G�jz�L�4����;�5��ϣ'?���@�.��՛~�l�����I)���d\l��Ѝz2t0�\�̗r�����-�
,��T�~��Ng� ��_0�	���T:������-����ͣ����B�/�bR��8��3�L�l�НFH��քO��?G
��2�D��Kho����BB���S8���v�7$��9h����� t�����:2e�*�R��+��<vO��#wӳ����`���Q���ҸU��ʏ��Y���z�y��f�B:>��l8�;��|����`�*��jVU���$md�����ò}��"1�T��w>�EnA�^�������.��yA��<1+��:F3r�nv��EZ�y{��ޔ���,7D��|+d�jtm����S(8��Ʉc���͐�O�x�R�c�����	m��(L�5e=�7:3��ݨ(���ϟ�>����.�8�j�9;5�+~��i�8}3�r!|��~\]=��J�ֿ��*>��S�F��jZ�f�O��o�Vܦw]�+�=oI1����'��N1���	LAmc�+�u��->%.ΑSǨ<d���I�y'S��]^og{$��p��ogI�B�ݽ[�F�����mŀpN�$+���g��RV�?��H֯d���m��#�َ;LI�_��в���+ٚ��B�R�|�`��Q�V�������e���I.�"�t�($�9�(�C9��n��N`���E�	�`�Yw1�����������ҵΛ2�I�cH�I��ND�t�����Z���O�J��� TъVY���T�!&Jp�z�����������Ú�}X�]&<��'y�6�����x.��v��~�A'����Mыa��Gv�l-8���&5�޶�%�Ȩ[8��7ramZ��N�/7��Pc��6Y�Sa�\RBȷ|S@W��p�,v`�+���~ ��ޞV\��I9�`x���}X.&Z{w���H��$!����jZs� ~apXD�7r��<tP�V�-�G�$�}C��e.��֗莩Xݭjs(��}r���v�fR7��z:{�	ғ��F����I<�J:B/�<���\~�!�j�:�]�f�}����f;Կ"�~���G�N���P+ �N�D��0�7�|/�t�[�r@gr\㽠4���u?c�0�ӷ��b>UckN��$�x��	"_u}ԓ��3q9wqd���5��%SR�c�w�mM��+备� ˛�AUn;[h���ɒ
_퓕�*X�K�J����/ޮJ�Q�zl��[F-|";}F6���M��G@�W;���Y<�{���P�t�/�ֽ/wa���W��ˎ�m��{%�yM��y�񨴁�����`�V����޹��¢�0�l�C�@�sl:�Vy�ekPa��c�4Y#�1+˝�g�JM��͸
w�{w%F�<HA+����|�SI7j����k�,@�tM#��ȏȧ��	K��N�"wO2�|��k���p�R���,�T�]�+6��
�����P}Lt�T��bVB�VK���{� �,W��:�R�#���oU�]��|��c-���
�B9و����~�h#�X�?+�q�o��ͯ�ϝݞ�����"tD����1T!��;�(���|�r����S�C�Z�P����bߘS����&]���`�������%Z���A�G`8ț�A.���t�I��q}P?�}"g15��ܘ�6T��З����TE���h�5u4{ �h9mWC)�.J�@��a�Ӄ��}��<�D�Q��kq�*��MIj�5Yd �{��b���2�ˎ;��BA�u���n�%�7��2ͦ�Z��)'B~	7�$�e)����j���uZ���W���x��`��d�}Qag��?�}`�:�%��y`���N���զF�Qj XBK�C����N�0��0cC �D�LQ�3���T��lA;L�\V��|��Ŕ�	���(���_h�څ��[����jr���7m�t�X
�@C���F�!����笠�
���}Zʹ���3/�|��������f�ף�|��A`u����W.�<���&�"L>{������v8t���+6� ���2B*��װC�^}��Wœ����F��je���Sr�a{`�����fѢ����"]Q0~��+u�1S�6�ԣ�i�no�u�cC���t�J�@Z=�,�kܦH���?F���v{�'2�M)K`@A��f���}�H������t��h� ayJ}:��*K����\�E�}X���v�=Zk%���. �����|t`�U�m�R�c�?�6k8Z��",S�T�V�Ŝ���ea���ح���Aj��L7������&����^�:S�d��e{Zҍ��\��Z�9׆�XJH�X�c�B%��S��r��8�ԼUT_��V��C,��b�ȍ��b{s�(D&���TQ��A�U�۶3��r�ȟ�#��y��W*�݅@���r
�$�W�;]�Q�o�)�< )�CAf7)\�	p���CB��x�x�e*��Dk!�ӱ�� ��n<��ĺ���;�c�ʡ���+FP{ݎ�������D�&��-�r>5���=?�:�q�.?���iZ:���F��X�|v��i�4G��+=��/�}s�x���w%hEL�@�
;�Mz=������@N�7U�;��[��Kh3珕$g���.���r���Tb�!�p�D����I��>���ﱠ��W�0("`*����9�O�֡�"�ϝ��6�+�E��8Y\aA]��84�W1X�>����.����P��%+�� #�j�����Y��X�՜��|���6�-��H��c9��׮(Pc~��(�����p�����0A�&��R��0Û8up���n���l���8�C���m���1�����L)�嘌v�q6�b�\�$z��YOX��S�.5$�Vr��Z���P�1�s+���2��R*^O�a�dԿ7G\$�N~�\��h� [׀�5�fll�t}GF+��x-��u��fc+���=Z=S��@�f��V�Ǉ���s�`�,�!�-�/��|O`�n����?f8�AB`�P2�+�I4�E�e_*���s�I2�Sv}-�ܜ�������UZ�l��KB�	�	eфp�o��{;���w����Addj�*��f�!�V�*��r��8�i���II�|�LճR ���=��{��2��z��b��ݧ�ϩj�)�_9P+�2���HLŞ�b�z��q�������,%�y�+_�Ȁe=����."��C����VY� "?��x�.��m��᠑���3��F�[4F99�;o�[+�Q�`��U��ө�y �{�� ф��;S�f=:�������:�ߓ����4^td�k�Np3��@�!��;�lC��p[�����obVj��]���22@���SM�����a$SQ�9ޕѕ(q���7��#��ݖ��N���mqBm!�r3�l�~��=	�9���l���vN���2��(%]~����\N*п7��h��ᖪ�6!Oy��1=}��Tn�
�A'����@��'Dɲ�`xw#�ڳ�5��{Mh�@�:�eR�1�`�V*b���
��KҽS��t�}�̖�2|����aSgM�f��[�m�p�������@��J���^SYq9M�@�H�k�N�}��lt�MM=k�v�����L��~��D�EQ~�3tH���6ޣyA�5��"���9�x��=���x8�s'�ŷ��f��>�W�1*4`�譖���ӏ>]�I�����2�?<�I��{φ8�o�9V��� d~Dg`��_��u�G�E87��_pS��B�����l;^�-��3Ij(s�����y	����(��@�w�g���UpT��y�v�B�>:7�	��0$�;�S���x��;l���|
�����YfT�gb<Z�S˾̦(����4Pv��8,�r��zƆ�-SQ�{«'z ���#'��9����5f��pii<'+h�J("�h�E$2�Z�)�d��;�n@ɫ��.OU�V&+�yw,K��J�.�R�2*ݫ�Vrb�0���Y��\���ܝ6{A����|(�8 ʯi�$��d�ϻ.�t*�����$-+��:A/�Q����ϣ*Px�2ğ��V3�Z��W�qR��&������~�,�J��^���բ��ߵ������0��n�t>[Ai���Ri�J�Z�c:�$�md��D�l^�^�?31#����it.@�b(5�c}�A�C�z7 S�6(Σ�-�.�yIL�$�6\���ʇ�ChΤ�\b��+�čgBM;��p��?�^�Ŀ��<[A�T����*����0����( ��)M���F���w! Q�O ��y`y�4V~�?��	�Q�	�2J�t�uI3)0�MQ�T���3���N�RܿyϞbwM�\k�hz	â�Y��j�Egf�i�չ�h�O"�䇠w��T���u��_���F�~�,�@��*j ��s0Z��O$Qs�<g��m+]�p�&YU�ϝ��]�`)���E�o�5��h�\��mW�_k/�#S�F��.+��eK����*��)j�@qk�h�Z\V��U�;�r��J�_�6=�P����/N
#��s!XKz�tVA�a['�n�)����LA9�RM��)��^!���S��_��>`H�5q���a9]��#@|%ϵ@�W�T7^�kM��O��(���[͕�T���.C�����/c@�����n7��ʺ��_E�z0�-;���*	Ep��3��b�-ZZ&��kw�fݫ5��ƃ���l�3O���N7t��}��6,��@8k�=��RpyW(���ݛm����B�,G�s+����l>�-������5��`@Am�%	^�(Q2��M&��o���|*G�Z�aI��(�I)RnGKNFi�0��/b����.��S'W�-�)x4h���q,��Y\y4JF�bOYia¸3�A�b���w�%����H��s�� Pm��Yv[�4��(�]} ��>6W:���F' Ӡ�t;��Rx�2�v�0�L��g�]P���.�w�5�^������c�h"��1n�D��X����v@r�B�C�R�+��(ko#ل��sĆ���u|
Y��P�]B�ꐮ�Z����=����W�-�_◷��a���v�SInu����šZWp�<�S2L1E9 ���ׁ*v�ZG�f���즳d2��E*8�{h(E�^�@�pq�����5���/�B�e8�=�'�{p�^̠�c�Cn���l%�6��P�|������:�E���|���)��gb�f8w't2���ڣA�	AE=,�O۸L�Og��%��87t:�^J��n�O���>-�w��D���*�]�Z�S��26	j~������.�K�t�ם{x��Ѡ���T�͝rZ�q�GW\~��o4�+B�JP�v�o�R{T�cZ�`N�[��8Ԩ��^Dd)A�\�}%�.�@0M����4���+�I��e���Ν�G~q2���(����g�hf���O�q^� �:��I6>�򨂈}<��|�jH����Ha�!��ɛA���=$�
����@��0	M��� _����n�F�/� ���kK�|��b?DXĆ?���w��M�
�NJc�x;� I'8����%p�ř��.=��2�q�rر���'���4d
Q� �<U���������M~.d�6%~#�)�~���	���oS:N]M0�j1iD�%�6��h6�򅟙2N���6��\<�����d<v��&y;uΒw� ��V�����m�b`+�{��K�s1���O����TU��~�C�o*�b��́��d4��$�8�����$��"9�aL:J�z󟳿���Ap|k�@��)>�-Ц�!2��
�d%e�91F���P��+��e3��W����Rʙ勄�澬r��92�m]��c��b3
���j����<	�%U���]j6�ձ�X@�/co�}8T�ֆ��|;U��B�e@ʭžY�|��G�;�/��
�������P�����U"���lSȺǊڑ��
#UY_�k������٨O�P�Pi0U�gi]�fҚ�K���zT��[D�x��4�F#��Y��P=A'u�����L��>����M�&d�<�����\�]Di�����S8����|D^wQ@�j��ހUf4�!��Z�N�X6u���oF�=�����e�������R\]��>�q��N`'�l�.��m�W�u���x˾�v
N�wi �EZc�017~����Uᣔ_�bR:*�D	�bB���Z-6�0N,G󉄨�1gy2
���Ч�{�V��stoO�>��L��at��4�����X�[ˤ�?�cUF�_9�SFA5�`(|W��Zm��'v�}x��+DL�� �N8[����&My�����7��MG]�\���Y�K�ز*��K�Je�D�5^��1)�j�����ٛ��Ľq��&�_[
���$x"�Ղ�M����:;�K��G*�9��C�q
�7!�FU���fHu�y��Zyu�u��R+��;�-�#'��
3w
���Xϸ��e5�'��{���D�F<����+3m���`O彿�>Ut�ql�Xo�V�����L{`WPq�n��"�u�@�k���1�׭�	J ��Uo� ,T4p뽏�D���	��f�\�[91�.Ϫ�0ڋ<R�|��a��v���	�J�iE��U��__��+��f+�#h4���^�\�z�Bx�����s�`��S�r!�@�#ۈ9kP�*ށF�W
s�y�?�:��)�����$�L��'��|p���~�$��>�C&�v3 ��q�� &���54"�3��o�����vΐ�*��>��Jd(Wۜʢ��A�⽿�:�L���H���?�Y��^0 ��Ά%��[D�ZWM�
�h��͌$�͌|*��~�!?}���{��Z�p1��A�һ�3�Sk_�������B�F�ˇy㻙����f�V����(�/�!�ʧh���X�)�f��/ͅE���	f�)��f�@fjǷ�*��J��3�<�����O��#�/7 y�#f��x�
=���ْ��ޘ�ׅ9��泷���(.�+�v3���U��Xn���q��|=Qn�Yy�քɔ������L���-s3 �7���K��;����~HyOJ�0��o&c�����SeT�pNi�GNQ`?a���e���k=�kN���0[g�}�~g"j�i]�9���Ы]����z�}�{���L���g��<�3��L3����H���D�"����N�c`q�$�cֽ�ݛ*�}�V���"�H��+z��X�
���]�Sd���v�+�� lU|Lw�������%��à��>*m��{��>��(�>x��չ��Y�I.�0��y�3�5R�56k/��K�66`K�r������D����t�l�e%`�B�N&�F�t�5��(��v�ڎk�td���U�_�	�rx��^�U�T�I�j��l5�Xt�ҋ�Emo��'�ݬӊ����(�P2ݑl=�y��]�Al�+�t ��LT������o<v"[�S�i�IY`9�=3�~� �0�H��ն����_�C�kW�<��q� �,&��x��'3�����v��]i>,�!��+r�R3haT�݂.C��݃��qЛ��W�̯����&Z�\h���},k*C�E�\�#������r^��AC}V!�o6'��Lh��"#���,���J`�b��se�ŗ/%���b�^7�0R�lw����NA҆��C軘ąYR�0��h��u�)�q�]����	? `�>���F����`S
Ý�9��D�Bf�p���!�nRɐ$jP�k#� w{��iJf�����Z�Z���'H�Lpa3w��ۚ1��c�gW=R�`Χz��c'�D�];��p>���i&�ʔ��x���O~�X��Y�U�����ɤ���-c����#�RB0��Y��;U/꾊Eo��j��{-�кc8�@�[}�=^t�pJf-	�SZ5)��1��W$�Ov�ҩ�?]ُ��ݴS�	W�gK':(.�[x�Q�����v>�j��l��m|>2p��>�d��e���h|�8krE6+UQW���-�>}��/.���F�"`�b,�Fu�C1�rU�}.�F�N�}����r�#���1 :M��٨�G� �CUtu�ve�|�J֋y҂j��k���S&i�`���s���mSI�SC�B������0Ug�ʆ�R����ny��(4��9vOm�MFtc�`��o��BR)i��:�����:����3yO:����R�
�V h8nz�EjiN{p垖�_����:� ���n��Lˇ"�(K���	��y�"+_���euH/�	;'���X1�<�b���O���,P�1����3��[�����K����W2q�e�e�����X���D^�,;2�5H7Hԟ�S��]�C<��P	���MȽ��Z��n8q���U���vS�fi�<U�?K9�|������>�X�����)�T�t5�����=��9����JN���\��-��/�r�K�ސ�-r&x@D@�F/	M���$���ĵ�e9���A�gbL��/l��,�"�Al��U��I�������oor5�u��29N7��]�Ywo�}��&���K�����c�m%�_ݤ��=2����������~�hq���r���Ť�y�úQ*!z�)DR�X����#�6}}��2CW0b���;&7{`�8Y��=&I�.d�yG�YL��|;�arD�:E��+H�>��Ο�
4�L�f����,�b��*�'g�<'E\��������r2�.���l���D�'&��~�Bn�Cv�����Hh�pr�k}��ߺ<	�9U���
z�WP
=�'Y���*�:���?�%H���l.(�ހ��.����+?uS��vH@��@��ҧ��R"������g����]O�B^/d����A	H������[����Lmغ�H"$�v|�o˰9r�#T�.�7!%/站e�1��*#5in}�p�=�`Y�急m	<������Tȩh$`\�E���y�B���3�e���'�tu؁�_�At����E�!J��*���f@�-�l�+
ₓ��>q~6�totw@w=�t�9K<U�A]8�"�DO�Vt�9�5o��Ƨ�d��ߕ��x,0���c�$D(���ݼ��Q��O������&7i���e6���j�Y/��V�aWʎ��Fg8�Q�%��g�j��M(�����A>h� n��.,mNx�`�߫t�g�uY`�b��޽�R,���%����ET,���aWf���,�2��1#B�36�~�:`��y�3d=���W��M��@_<���R����6.'�˫��D�B������R���̇0[�=�.Q�1�)�)>�H�^�Z���1;�$vo�iy�b�]�>����Ff�f�Y�C=�@hF\}��߯W���ky�N�SGR���#Xa��seB!R�?��o�k!��?gixV�w�1u���L�U]�����Zg%���ss.D}�c�o�����xZv�]�2G��%U�v��]8<2��>����1����4��ǖ��,%J��W�V
�iU�P��h�>�3�/���U��Hw�X����sQ�A��N?���jqM�PIN ]��U����,�jXq' ���ؓ�V��D���*f5*5�x��i-��CZ��w�@�y��7Q3�!L��٥��u:�A�Գ	���K8�����Ħ���aǰ1=�#O�����6������h�C�n� ��o n�]�셕�f!KBG[�c�)���Y/^G$�H��SW��MF�!L]�^r���MO	��������Mu����6X��q��m/�|?����`�Yj��IG�p���`AN�ri���\gITt,���u�<���ֺ
���{.��%-���%�/�U�����a,��� �Tt�����~� =CB
�il=�b`3.u�!{�zHY����C]�2�#`�9��Hf"�k��%�ÿD7�?%a�K��5�V�r��j��k�z���ڽ\L���>�y��3�j��~Ͼ�.���D�Z���6[�e�;(e�;ң�������랴O�b��f�*���I%��x��N#b����R.8AA�S}t�TX�{�f\}x�'\*�*������6X��w�GO6v�Z}V���<2J���Ϻ7�t��ؘ}� W��ҙ �K��; �#����ȖОP漋����q��2��62D���Q͔�'����eٺ�N���Z�ob�k��^��ov#Vs=&Ά�qmE�d�4q�3?�5���Y��N"��f�_ν-_˿�<[�G��
H��y�}�J�>x\Wm�ɪ@�%HF�br"ő^�L�Sq�Qy�WY��6���a3�},xN^����kW�ߞ��p7�@��*Ҹ
�I�]<#hc�[�C�ҍ�@�]��(d����n���$4�Y~t5��ﻈV��adah\���S9k#^nՇH�a��Ue�ׁ�B�,�d�8lxx�_H����m�X�1ߥ.+�xZP�J~���<n.�NI���^ ��F��oPA��}�4P�r�2I��h���J�`�4��� Da!K�`h��n|Γ�)�%��*$�HK <�6��;z�׿���*sl��e�~�,[�3<�5��r���hm+�V�;Y���?�_�Ł�ٵ6�ݍ�B�8�q����V���|��Hl\��
"�C�?p�Z�I��PA�C�S�����!E���K
�����A�I\�!OH��J��=({0�J|HM7��+Գ�W��h�03L�>Ѻ�Q9��Qy�sM�ގ�ũ��5
 ���=uI�/V7�Ʉt�#~`�Z����jH1|�n���d|�ۍ�T�6�M��v���c4�K�1�O)�vp�J����{>��3s�^z�3v�� �gܔ�nF#t_�����.�քR�06�����M6Q�	�5򣍁шr����}bBf8<a�h=r����_lW�қ~n�W*[�/"����f+t�j��GGR�q�����7�V5�2�wB9�r�4ڳ.,D��N�
�q���>�ȞH�끧0�UG��Ǖ��(М���ޓ�@+VRJ�+(�Y��}-�޺]�BR�W˳�'�U7_a�&��xp_�����x�DѧF���`yuI3� ď�8K���ݣ���M�T�:x�z�r���亯�:�U�`N�0���[Ս�QH���ܰ
�h@-]�Ȉ�C�i��M)�Cm�a6c��w�v��Je��aC3Msẋ��B�He�t�{7n�a�� ׭AoL�Ɗ�1Y��r�4��hƛ�G��4R�*��FR�%[}W��${-q=Df���z���~��j��*��B�{9i�:����P��\�$zAsT��̅���@�����%�E�k��3aC��	�����G{n���Ù0[�����s��
����W�#ѥ0d�ПM��V��^�K
s0�pl���Jj�"^�9��h�;u|p����m�T�F�O�0��o"��Ǌ?��T��E v��R��zn|>h�]}WP�U,��1��ĝO�E̳�`���AK�d�[���3
5�YX-��� �._����),���(�!A"��=�g�����8�d���#4������Ǯ��#M���"�����ԩH��`�}�|��ّ��S6��\�W���+�a�}¦h�R��Tt��ph���p��9R�g���n�I�ejxs�E�	�L�f^��d;�6b݋ܔx�e�a�����~e�%��KC���������n��&�|�Ά>i��@��&��y�������
V�8qj�ݿ
H=�����7�ϓ���^U�|I�v*��yO������7�&f�\��8��됚Km���g>�]��S���I� ��x ?���(��F�H�
��F�SRAEΊ��j����	J�*_7� b��14�v1�k���z-��̝U�~"�m;T��e�Y5#�wKrMS�h�?Q�1[��N��"D��nQ�����hO�ր�yc;�l;b�)=én@�ŗ���$tڠ9W���!�"�e��i[k��f�{T4�d+&���@Nz<�VR��/��4Kkl��:w��g��S�r�|g��1�L�w����[8#|���hRg������dǔ�O]bP͚"�W8�O}r靀f�����?)@��N�fg�"�f;:8Յ�U���g���qr��<�6}�Ѕ����#�\��+~�omO�z#UhjE�����̮���u$<����w.f4��֋����^W�]��q���m,��0��0�ʶ�#��[k�0;������a�p�g�0�����Z;Loy�%چ}M^S�z{�+�{�:�b��ѕG�\k�o�	�#�����������R��.�&MdU�p�"r���I�O�NumB^�qm���X�Gn_�i2,��r�͞QLn_ ��2���t+��#��H#��,��Z ���Nu�I�s��w�]	U�)X<9X,��k�%��֌"�#���5c8��o�ՠ�C3d�K����)= ��}TZZW�˧�l����v{-����H�h��@���W�VPs�!2���~\�Ć�A���q�Z�j����g�BNt�AN��ʊ��E~��>��\��Ef�f���Js�i
f@�W��qޓ� 
���`��f�ڟ�`�p�K�t�$�JP_�{���=Fqy����Ls��}M���K���]KTSt�m$u'[n�#���̫��G���+\l3��f�5�T��*��]�x���#��xLC9�2���2���T���ZK	]�P������:yp��b��C�c��!��X��=?wt��F3���F5 ��u5����η6SP[�2��L����ʌ��҆�c�Aoʋ����+4�� ��;_rB달S»� ��ݥ8��S�9�ö񎯱�)HW\�dzIx�Do���������t��ɍ��&��VHc��1�l�8z��$����f����4҈��^��Q+<;�Ѫ�>@}6��Km�8w�D�&D´f�&ш�"�G��!��o�vxܙ.�����9z*-��:�gs-��� p��*�z�h
>>� M�{��j�i������nh"L�
-��C����Q}=�|�n!:�V۽n�wz-�Q�'�s��7��;Ó��آ�����=$z#"����K�@�o|�T�2'�	d�Y�a�����\v�œ�1������1t��}ȏ��\��'��o�P���=�I2��8Q�.?j���l#9�S]�2��6��6�C@ ��3
M��4����u�}��ܡ��:�֔���*!*�L&���
@���H*��H���M����_g�|IxmmG���b�h�G�G�2L�!�  �Q�~ۅ�W���'};tZ�*�(��U춧r�� �]��PW�y4S��٦�0����L��m
���Ho<�b��'��C߫�.Dz�N�>f"�D�j`�Ď!r��P��֢��ż�@�gahެ�#��+pc��y-e1��Vqy�KJ��9h�M��o��p����{�I\z��=�G�2r�Y�ΤT��l�
8Jk쎀P�����.��y���`d�Ӡ��r�)��7PZ�d������\�D{��5��g�Hp�z<5�?d�oK����i`�s
���"�|^~��QGR ��<�L-+Ɍ���hu3s�E��n��Yzt7�Q�h��yR�H��N �CZTE��k������G�5$/�=dM�B�+������?S㦝rXĮ4q�Zȶm�^��A�5A����{�ݪi��r@�9��ڄ�VMK�:|�SN�3?�XT4���s�]R?�x�E(�8�����Gۤ�+L�\�5�G�=�<'���4�2�(�Y��B�6���0���iz=�`�h*�����Q��̝��O�j�{���vg�{��e"\�15Q��8���\��<�N&����u�FZ ��J��H�xk\(�n$IѥV���ra�l?(�Gg�hO�3)��!I��f��Q���Օn�Sm�J�qhT#U/U���(���_-���,��b`U-8(�9G�&�3��ʚx�hš<V��nNi�Xi����o�����`�f�1�H*l����'U=��%uc}*��'n��}�W�<��GDP��_��V֒wPlAnG�5���A8��_��=��Ѯݡ�HjҼ�l.b�Y��������*��J��-j�.�zv휨ߒK҅Y��/e�6D�����j[S����i%[`���@2�ƪn\R�
�� �#�W�$�m}�I�=����D�M\M�P6{�$W=iR���D�"�V��lh�Pd;��{�]�����[�ߕd�K���$�5%�� ��I�"����Un�ۀv0C��|��93�%�X�i�~!�qL�g���`Ku�5�����J]."ﲿ��3�ˑK:(�qD�XΟt$#x��GE���SbQf`\�]^�l�
��z�vodw�`�P%��0�BD��:����
�[`&/��#��F`3�9'�����07�m
�ǵ٘Ӭ�ۍQ��.�@��ji$WPH#�R��3��\\{w(����d ۍ���h�#��X�,Ӻ�=�Pڕ������d�+E��F�Z=D:�)��r]w��bֆګb�^��㵊"LH���q��SюV�l��/����)�d4H����? 9F��]a܍�D�%�0ӾjՃ_�y 7����c���,森X�s2�����Rn�X^{�R�q�h�v�t5~WC�g��^i�畈'�[��X�*i2����g���!t	%xZ���M��pw$B0a�-�IH�	� hhKУ4�����<H�tջ��4nKH�iw]�݂q���$ӳ���D�{V��~��J����8���73H?=�H���.�u$�[9�&�e�o�
����n`�;���ah>lV%x� ��l�9�[d�+��#�3 ux����(�~����;DB�����;S��W�P�L��BM��Zv{i��tӝ��(��)�%�8�X�Q���<�3�: �l �	oC���3p���Y<�U��:Y]ə�]?�"YWX�v�^�o��pT�cև�YG}����i��-Æ]&�:Ag�3�/���������P\�Z�ob� ���c(�4H\L���$��r��i4��0��� ��ZԱ�s��=������Qyf%h~{xU1,��ս0#�HЎ��s oo��r���Q~҅d���8*v�
\��P4v�3O�n`Xr"	�G�Ғ�,���7�
��J�e����"[�R����	I7�b5�G���.3.B�NE��]dH���B�"Ůz�k%B�NS�x��*�3�I�ڜǕi��8�zg� �A}�9h�C~e�in���K3���W�e�����f&!7*@�*�N(3Q֎3, Zo��.�V�˰�,�՗FfE�1��ʓ��_3G�q͎���4V�y�����Ui���-�I������.'�Q	W��Bp�~$�Ĩ�ft��|�������pem����T��X(��7�����Y��R��h ����+��Xi��#�J��j^{�����E��|����7x,'�J�x�� ��-C�C1��L͑s�^�˗��ڲ��eѩ�v�X=Ɨ �2�E-���D��?��=���=(#3_m��*�5���@'��A�.BiH :�/�Ĳ���������H���eQ���8����l���JP M(l�s����TY梦����@�jf���9g�X�p̃�8UF(�ީ���$�j �|�%��Y�s�U)s��<7l��ӿ[���I~�������-D���ڃԳ�Q������ֲ3���HȞ��{'\��b����<�<
7� ��=�4�a�6;?�//�j�!%�6(���>P`x�sn)Q�G֕�hG���J��$��
�j�I ��P'�l�.�	�t
)�#��a���U���H�ζ���M��Bz�6�^X9L����B� l�HkĎ�i��dہ�ҙ�t�|W�D��~��y���Y�k���sY.I���a�C`etX:���{>��T5����p��6���P@�����R��a]�3�{�H�f��u
1W؁y��]m�M���ޛf!�{�,��k���I�z�5�M}�bG,��LX'6J�I�W�����9Iԛ�L���m�7��P���M�72�.�G+���v�<�n�Px�u�,���b�p>Sq���U���x;�,S@B��0g\���m�q^��eڬI����.C�diQ���{��l��K�"X��f��esl�}@LN����7pA���P��XЌ(�+@���M��{�b���]�1���;!3j5��}��_�Y4M����[�?�����C�zw;��'������&T�ry� p�\P!��q"����b�1)A���)؉h�[�M��Ͷ�^�SUV�@�,tW@?Ne!�l4J����l�!��^�V�X��R�x��E-�>l������x�w�"k���X[�W�dd��m���&�G�\; m"N�&�N&A��h^f��|L���pӼ>��{9�����	`m݅htV,9��J�'�%U��u��6�/ÂM5��ŠL�d�(5R��h��G�k��3�p���+���#TR4�i[~?`"�@�όT�l5f��2_r]�	ޮV0�c%�"L��-���&Iv�o+����OB�����܊����J�ዮ�%�|��7/J�+x3�K��38�q���ǅ�B���G���>3�E��TlO�~9ڍ�gĜה&om���"�D��
Ac���7b�(����߂?7Qg�t��r�ҟ2����ipY���[�t�d�0�Om49`p�X�Y��$"!�Sl����?� ��j�|Q�T��f�1� �V���J�����n,�Y�js_j��ws�;�V�͹�(!�cUSוּ�(�B��E���_�r̜c�՝��@�^C���EB^攄��mN��»�y�M���E���� ���Vtz��K�[����t~\F��:e�Լ��-�ѷ�=�2�a��Lk�kҼ�h�59�~YJ��H�f�Pk�:�$��"]�y����>nh�'v�p�o���JQ�Vy�g98��J�ó5H%�}|Z)M%K����d���"�rNK)S4`�ԗ,V�T�0����<���0.AL~S�^V�X�v��y����:zz�M�J4A8��Qʞ�H>�}�9�\�:g�v�r��WR�M끲�\$&E$Gw�546�	�"`�չ��]r&rz-?QT���ۏ�!�?w�Ư������!4�
�bj0��wձ>�:�����kJ*#���5��;T&�+~ɔqi�dA�9]'�����ت��i5�Ə��d�׎���|���| �W�1H0�A�	���]�B8EZƔ(�7ߠ�k�l�2"�dD�ZN��g1O�ۂe�]�F\�Z��pXK�ф�ᓩ�y�Z�϶F�C��ML��L�q���?+����5��5�~��<�
����	3��I��[M�`O��}HX��r'HIn��{`�u1�G4�/�����"w��@�d$B�������M�eF�{Xz�����WnF�#���{l�"�g�Fǯ9ͪ>E�,ݎ�J�C�Wҁ��_6
���n�5] ���"I)�r�BH�]6K��靛�{��8v�L�r���f	KG~�_�3���wꃋ	8���G~��r��z�`��WgP�.c�$�D��ǐ��d�xXZ����Rg��:B!��d�h�R�%�(�JZ]Q)�E���������(�X������c��b� ��r��A�]��<��!��g�z���|�gL4,'�_�Ħ
���3�O�zw6��N�,NY�_��; �YY�$�r�d����C��� �H�AJ�
1[�N��Q��O�?=�?<O>��os|ނ�89 ��C(D2<��2!�]�v�#C=03�xӘ���͢N� S��^�~�&�FoբIk��h���y�#��B���N���(�	 ��C�Wu�a*�$��L��Z��"� 6;5h��S�.�R�؆Cj����?��78ϯq���>�PNi�_��Mw�ՅF���-@����,T@��{i[���*��7���v+�-�3�e��$	%,�|$���_UY��ek65�&�3} ��M������� ���U��R��B!N�9����V�zR��ģw���L�$��`kO9���P�V�$�s?6+��Љ����\8�b2���v �i1�F~B�9}z� Z�Қ��8��ӰW��L�մa%���|1�a1����!���&r��%�ϡAg;����}eN��D,� ��Œ*����
�D�Qe�Tf&��������i_R�W�� v|/��P�����������,�y�̒z��h�M�ě���H�@r�dy/�,j�c�W4�߃��n�ߞ.����=�KΓ�Aw,��|������m�H$@]����'�@#y��/s�T��IoDzE�W$$���L�>HK�3x�2����Iyy鮳 ��_z�;u�����j��o����PJ!mL��
EtbQ� I!jX+�ko,���3O؛�7=o��<7�]ʴ	���z�� e0�X��mÈ)L���r#D��>�P�z? ����j9Z��k��ʇ3q�,`��5��b���[���� Ѷ�^�2���@F�������.��xtK�q.�6����j��Wg��Xc�-'��al�%&`��Ig鎢͍+n�<6�~S��|e͹�
�VE��������SdXIm�]�U�BzM#��Ya��'���M�^*^�W�	U�iInQ(�?pV�ƺ�UD4���&x`m�\����lsR���Uk��5֞���RB~�l��G|�Ҩ��k�ʛ��T&#�TU�5��!��6��/�D&zzA9�z�I�B�A)w��U"5Mһ���?؉x����.�ui�������A����|�*�F�����?>K}�Uo��ޡ���zS,�+�A:M�'ݣ�����rg��OBT��|����D�v�%��,"s����n�7�	NT/�qN���PH��X��0��r�r[(q����(�@��G��wy��-X�wprJzB�z�	dۯ+ٕ��ϴ��ǸĄy�+���J�;tN����j�m�����|�m��/�^:]���p�	��&+Їӟ^:Hs$l�3�Ҥ��[�p�!��	���H�3{����=i9��CS.�e:O�^/��Y(H��s���"_����0��(�RH(�1�QXS�֙Q�����~�$K~U��-,?%��x)�����:��?��=��j~3�dVdp��f ��r'�o�#�Y�&�<�F��R�
�u��:9�>��G��\�GR�&�9ɸ����Z�$^��铒)A�L��h�p�'�V���>r�Bqf{�0X��;�y���"�n�*w6֎�=���v��ܼ�f�V�2�e�sPUF�YbO��[���c,w��$`��o�,{/�#{c��.@��r����|����Q�<���Zz�r�
^�Nb$~�NǸo�
K{@XD�8��X˿sEML��5ѷ3����#�H���R�-���^#�Žḽ���P���Q�����Ҭ�ˡF'S���={�k/o/�E��g��qTA�9^E���d��u��`���a��zە�;�\"y�>7�ψ�V[�f lFMsrS�g����K�Z�㪅�.���!�u����ܟ4�,>G�ȯr�KQ�#z�u��+|�ζ}w{HM��I����W|� #��i*�B�*�B����l�Zl_�9���B����bܚ�m�!%�ڻ�j%�"�f��V��!�8Q�wd^�o~7�H�Lc�u�����:D�5�X�X�N� 9���;���%��$��LT��� >_W��V.֜~c�J��D����޼�����_����ݺ��m�Ge
�%�.>�Veѫ�?��2�����+ȅ�W7ײ�7���tf��FGlR�Ӈ�`�Qk�>�lڊ��$-/k
���'��H�v30��v�C������Ng�l��u�-g4&����ӚA��g��2�e���nX�N�mIC�X�$����!ѳj�V�i�K9�!1��;��8�՜�-��
�0��!DO��8t1?�H�z��t	���a�6�h���B�q�*I��9���U������Z@t��N���3�؂��|�x���T�\�]�������WZ}���ڌ���&\���s
�c��:��3�T2'������Ed7���&����
K.�lvF��qX0fټUX����+����heY�ϧ�;'Ŵ-%e�xP�u�Vd��2�A�C����f-lM(��н$��O�ֵ9�J�X4����'��3���ߤ6 �9����P���|��2�`���fw.8e�8	�\��D���+�i=3ɟ17J�&.<_d�����M��-v(����<6�׋�3{��g%޸P&,c�]O/�g�1J��Yd�>�Ge�!-c�H'���C���Zׇ�"���q;���3`&�Vؘ��C��N�6��BNhХ�C8��kR����iD(ط���O�� �~5��u�����nb5Z;����Q3S�x���%��A3 9UwFK��l��'����́3A��cQ�_8�]>�[� $�����ġ0< 5O��xB��u/-�M�
a�.��p�9~o�~��n�kD$�G!Oe.������*�N�n��+�_�P��j�p�7���h�s�˪uźȉ��(��R���O�@�Y hu��_��	&0�6�
ⴗK��[�zMn�N��	����4<*k�4P�s�*���-��W{�G��L�ˮ�T�׹V�RA�BŻ�RU@A��&��{�,
�~q"�\�ߺ�0q�l㙔�͇Ne �t�����+E�.���0(��(l����Q�Vu8K�����t�Z~�����	��6Z 7}%
[L$>��5^|��{�����SJ��B���v$~oUdX"Ɩ�b���Ä�g��g�&��i�蠤0إΰ��?�,�3,�QH�\�5|aY�>�o�fa�b#���"�D_%��$�ϥ�T/��v�2p�OL�|x�ul�nn��*!݈�8�7�-��,E��* �y��;��x=��⬅��<�M���0���䏀"���9�JQ�S�л3&�	��$0M3I�b���32�_6<��#���{X�����s��4J�b��4;�;> �$�ʓq-iZ�N��l')�yd"j�/w��)��էٓE�]�LQeʂ��4����rzп>`$�l4`)�G�pN�4���SN2u=�h�&�>�q&K-qic�Y���%f(M(�Ȳ�y��:3u(�\n[�2�S�ҹ���H��=o=���Ql�fm,	�A�MЃ|��΢5� /
�QF�[P4�0�o��?�}XdzA\�W���<�	:S��u��ˉ̥�a��E�bC���Fu��"����@�"Hh5{��CT<���m��5LZ�i��nv�$&Ћ�P8�?~Udz$�\H.�sjj4�J<�`C���	�<QIPCIp��n�x�c�J?��� ��@Ӓ\Y����-��W*���#���ن�U�ڽ�.�Cy���ٛSv	��9y�L�v���͑�]������#�A�0p] �"�̗�9�(�l,U��	��b�p�Ri:-�R'$��zU�@�Rܪ������1�;�n��µH�u_MXZ����]�Y��ќ?�d.��l�hX����#��^ݣd(a:��@��hT��=&�k�O]��%�u���<*�� /�pU�P�w���񚎞�M�U2�! ό�!nh�e���6�"�Y�xG�R&%�}^+.?��� �5�!��-\���rRG7�l7����xs�q�ׁ8Ed�PD\d��_]-d�^����9�����X` ��?���|��3��e���������4����[$1r>W����$ؓ��Y&��3]�;I@��'���ly�'!ߊ�i�Sn�ج�0�x|1��x����oz��B��\�=%�'m�+c���u�A�nbO��7}��g`^������Ŗp&�f�T���Gϛ�Rv:Q����I-Y
��&���X�~��h�)`��������N�3W[GӶ��T\���=�Wh5п$z��k��q2E��gŻT��v�����g� �N�W�g8d�l_/�7��x|��$2"o��2V��:8�����|��Q��"����p�N��A����j�خ��Pn�S��/�l7�#��𹰲-̸=_,C!��a��Dx�� ��s#�U�g�=p<%8�z����A�,}̲Z�j!�@����W����)�f7��|S,���|v���hcf���~Qk�HѸ��+�7�6M�-��h�0�zV}н�B�M���n�-��s���+�O���&m�	��>� �)f�%��8�.l�����c��m9�[b����7�3,���-�{�D�/��R�vx|Xb�x���cP�U�<�NivS.nU�� �).��U{M�6m��Oϧ�/4Bl�z#�o�f���Ob;M/%���r���cR�Ón�m���	�z�ۙ>�o;��S4�$[��ǚ��+R�N\�5�3 ��,y�J5��?��C"E�9�g��9��w�υ��&v�e�Ա�|
���1�=�wU��^�l��8�sbyd����?=-21�qVw�jt�E��Ybpp��`"�PיV~��pΑ$,$;��8��%�M7��/�wΗ�7V���DpY��_U��X#�����Yw՞�,���2�"R�n,�X�����xb����\�쳵-	�n�5�҈��n�u*�>rx>j��^�#����.4������^��m���o	����.��e����i�2Y&�ҵ�7�?����um��l%|�f��&8jd Dz���d�L�b.��a�dL�V+*^1�co�Ҋ���h�b�\(��븺�o�u�X�Z�	R�ԡ�g�T7��t��:�������?i`�;�amwج9�m������-9�4������e�����R���Cl��q�=F�6M�d�Aլ\�'�1�S7�h��g����d�[X�<����F�X'�������h�a.���g�E��#� ����:]֙��e`L��(�=Tt�Ϥ�)���m��G�	;ݣ����M�VI�ط�2J��z���}kɼ��wf!�N)� �SdZ��}�n�`��M��K��o�+o�P�殀�1S�I�	��]�?��\���6�4��%��Yz���X(���f���LF�l��W��4��y�FSP�l������E���$o�	A�ŷ��/|\�|L"Q}��L��Nm���	�2�K.��9�E!V�J4��VX �va���A��Ԅ�2^�\T�M-/��](~���d!B���\��ug�I�JdԎ>�)��N�pxzĨE(�}�TN�F���� 2}b�3?�P4�K���2�X��^.�"b;]�h<��x�>!)i>-�뽾G7��c:f{��M�[�������x�.ZF5v@0�CS�ʭ^9�~��H���YE����W�V�XX5\�&9�����#h���h�}�P^��e��b�gp��?,�w���|l��2Ϧ�Ӿ8'nUǱk� �Zi��^��T?�[��rd:TADns��j/zVy��G�+�L�7
�����R�W���;��!�+b|��^o ���ҝ��/��B�~�c���g��< ��i�CV5Oc�i��Ֆ:Cz��|fۖS6�0�3�x`����+��>�$�JH~�O�u�}FDq*��~��c}����dJ��B�� ��&PrH��ڎ�l�"!�)��b7����$�sv �Z����dp��q�[��Cҩ�y��G�})����*&�تS?#p���$�j�$��!��v��W.����,�?�����s������lU(���q���O�e����n���/`z�TW�0�*r���bw��F��P��	��纖��$$���u���"�Wj2�������� �Y��ڬ��k�,��:H�~l�v1P3��R��
�q2����@�浯/��T.��c�=;��f�!W�^<�����t� 	e,���hWt�)'�2�_�p%9��hT�َ��GŇ�W�&"S�a_�>Uݙ�y�<�뭚Q�9�R}��e�Յ%p]��1��l��U(ܮڗW�^'(8��>��Eی��AcD�u�(0 �Ӟ%=��7s��(�A����B � Vϛ��hȭ\tuqt-�.q YS�SW���.�����q7H_$=H;����۩��q�[�(� �f1����V�۠�4�Цusk�p�{�<�Vb>FB��'6��1ц�F�[U��_9��܁�ҜL���.X�О@�{�@��qV+�aĄ���q��lu��<<�W4�ȝ!�q%�u������ѺMwI���І��0sb��t�F�oE��X;0%�ʵ7�-	�jb�DI#��A��R���l\�HV��dE;�ӿq�����z��5[��Ԃ�	,&��4�"�7���˫�:�͈���OB��� N��<P�&�����~a�٨RP��l��T���R�{���|�Ӊqg���*��NDsR�q5�8"6�i�Ě�	B���)��5�pL��� =+��C�7�G`�*Ҏ��9�{�!9C���}�~n�,��|��f�]�Qj�
���#���+�2�Ra�!PJ�m������]:2�����U�Li~�,���C�e�v�:vA8q�ފ�Ҝ�Fq�Ľ<v�)U ��� ����y��gu�A5w�1ޓ��:�O���Yr���IxO�#/ɈV�}��
�W>io�1�%xx��/�>[�v��v�@�W\P�p�I;MytX8�2��d/�$Tޅ�f�x�n�{R��и��B��R �R?(�I��N|�S;G\�RG3��R�O������,��$gs�5z�\v��MD�=���k0�;Ґ̰S;�£ک`}v v@R�!&�bڰe�C�i9i�R�9��w�sk%g�|����ȕz�R�"�
b3�ŒoL5�d&�~ٻ�{��BF�����l!_�MK�'h���E�#�ҧ�88N/r�p�b�Ȳ]D��/$��,G�<�ё��=B�6G4/�����Y��e)t8ӹ� �F��%;;H�Z1:9�W��Y���U��n/ajrd��
��Z�d���G���h�Il�L]��}�{+����c�w��ZF����u�*P����9Į��. ?
^�`̚�y��E����R�x.Q��	}�e�:#��z;�^}
@��
� %�y��9�\�����^��}J~��1|gI�OK�ը��n��v9����bgB{]�!�dO�&S �&����+S�4���7�+J��w�a�ö4�'�~,�gU-M��k�5J	���)pt/�Q�h;�GG��`���$l�
 'J��(��	��V�(��m�p�/u���ؗvc�u�i3-��*��(��)�uŖuj.z<x�p�/�p`����S�\qa���r{��џ{����bTj�����lA͈b���#�)D�9@��x�p��|��6+U˾�ϵ�$8�?��Yo���?�8r�2�JUX�j������&�U�[6s�<��t"H�8)n��.C�����4����2eMiayu�-e�	 �vg6�=d\t�ݭ�T�.�ę��_	�}�Γਂz!7bfMד_s$�V�7w��rgQw�};�h�虚�R�1�M.��夋`j4�b�P\*\���|Q�9���x����}��Qs��Ok��@� �{E���Kl��_��Z��d��4���;m'�@*�{���Տ 1��ݰ����O��D4�t<�7�#T�t���Rk�@hH���d�I��}�X��0����@)pk����TN�	��1��]g*"��i�*�G1 x��箚&P\*��\
�k~�h���-1�[u���)@>�+&�s�(�+ ��*�_?�þ�@f9�㰸�ȕ@�x͚%B��DR�
)[��T����K�O�!�t�M��ΎXO����Tͷ�BD^"Eb�l1㶣��iG��,S��DP��0����c�����y�6�z�Q�W�n���l �1�`�y/��7L�χI�	;��!�����"x��*ˍ�����}ދ2h��W�LΏwF�ɀ�^��6�s�0���X�昌2�QO�I\k���	b�d�_YEުZ
6�l��\8Y\��J;�QU������R���SOcp��Xm�h��q>0��o�Z����fyq+�%����C_��o�v�o�@�0W%��S�f�> �(���oF����Lч�Z�]����6�j���I�`��,+;+��Z^�#}������h���\߸V�n�/\�`��|���0*�%0���|JN����W&H�z lI�G��_��k�v����R�-�܉{J>�h?O���4^�t�+�����c��V+�������ވ��I8%W�h!�'�pg?JX̴�[����s[U	 ��M���e9
M,oW�����ϗ��d'p�UK���xU����7��|�<��69y��+�I�B��SQ3�Q�i݂�Pd�P�/�Tn�Џ]����c�	�',��y�J�M�-9lK+�oh�0���Hk}@%���H�2E��?��.^ x� J~4ĽJ�,�����'�Q�cB�C�bY	���ؽ�_)6��&� ����.��"g�
�ǫF��[��4�������J�>�@����A��A�Jt@�9ȯD+Fi�nΌ)���o���)p�F��%C�ࠋ�I-�1�8���4!��]�	S�f)Ei�3�z+y<�2�8����T��N�����tN�a��K:5��/�a��YB%W�1�y,���}Q��b���6RxtR��h�BD3����1Wp���v����t�h�`�~�˯��u����k�Ew�F?-M����kPV���h�f����/�[g����܆��>�0!����(�Y��@K?�0�ȣ���_gf21'�u�R����~���8�(~=�O��e�d�?��W3�R����.a*R)��OU��g�]�G���yBC���g�q���mS/�ȫƾ��[|��AE�ZϼU�sC/ ��r�4�ħ�Г�ñd=�QOM+�&��aϣ��J2�|(�r���<�7��3_G�͜�Hq�v��;S^ 5�i�$�~�Npx����z/2<���q��芥�5<k�~Ir�C_�����]�<E���&=x %�{��V� �����?t}�����cwPt$�UvN����e$�յ�K#�K7D��:�/(R��l�	�������i䒄�d�=��
�x�ʴ$a������ċΈY$К�D�E: ��fF.'��_�x���n���j��Ǒʯ �!�Y����׍��D	�vgR�0�)�����a�Ά)!O�(�U��s�X��}�c}a�>6�:��G���<P>^�B�Y�.q���O:`~_r�Q�T�#C��W~x�xK7�ټ5|]D65�rL��u�<�E�N�0�: �~�����ۙD�b�L֩��x%�,��'�ΰi�Y�կ�T$� |
�TR�O>ǀ�/�q��6&y
�Z�`Mԕ0�+�c(tDM����=x��;3G��0��Eq�k>��ʧ�Ih��f�uM�t6
���Y%H�F�}�cC�p���d��	�;FI���F�Z��s�G����m��4T	h�wV��o�	p�£'@��Qy���C��J9n����mh\�/��פ�eT)��()RF#I�����$��sc?=���K�����v�0��'�o�~�Jt6�o����p�X�����@��l4�7ew��t@<���B}�<�F�y��qY8�g ~S9���jq\�a���"�p�7�htU�ޘ�6@�)X�1D�
�gB�+�GA-�-��{-�d��w�iԢb��h�"/Rϛߢ�mK��BF>F3w�B�9Mk޹�����f���x�'p��N�W�-f3�o�q~B>=%���������:A���s����g�*���7]�!�o6�����ۙ���u��=�����(u����|	Z�U�ð��a�A_>$��@�QSB�Հ��X9%{�Dë���d�j*+��i�Zl��;7Aje,ٱ�A�E���¡��-�+�8.����4�Z�L�7? ��M�7�n@���3$����{�P�BI���e��Ҹ���6����{�Al9�l51�wl6Mf?Od��yǪ���e�o���`�K��S�l��Y���	�u����}��.p@�� ,��E]گ�e��@�Nl�:(<�U�0rɃ]��G/�%2��'ɋ���m��^"�xS�-��]�_��A�ײ���0A�}gt���Б18�?�`=y�t�sG>�b[�^��}K�Ƹ?�~��v6sr��>J-����4�C���o:��&J9u��}��x�J���C�>6��t��4��@_�G��˽B����\3��iŚ&���h�{���M?B5�v�'EhV���[c4#�� ��G��������[��-�*�u�Fz�#�������Ӽ<����V�^�������n ����'�C�iY#�C�B̖Kv�PpI|�W�aK1C<���c�|A�Q����+�������SD		d�[�[��! �1m��0
�Yf�C�L؅��gո��ELh6��h}a'9�����G�i���t�̙iWKJ�g�BP�!N��W��fiJ6���+F�Ǯ���S;w�%��*�������\Sy;��c�Ok������fl���5���::9���YJ��j�٘}�{�4����3	3�O��?6���~�#N�fh��������<���T��P�29�K���JP2�����p���܏���Ss�H�K+-� 5�����*M�?��[bѐj��J�"��!S}z,�hoR���������f��ȭ=`�����?RS�ޅ���a��$���9�����~�.cF 2�����gۣJ�u�hKJ��BρWQW�wd�E�"�$�����]c�����4o��u�K�hj4���ߺ��R���^!���G�,�o��
�P4.�ZE{��;�C���I� sK/f�2]��&�v�Ys�������4�-����eʱjE�!~�c�<��܆~�0�����!R��'Y	U/AB�*u��d����j{	�'��C��]ȟ�RpR�	v������n��ƿ�!	b��]��.�% ��O ݴײ��|	����@��$Ћ�<���p� ���}���Y�h�QJ�֤G^lw��GOR�4t�˄D��3�d�β]�Әe�Iz..�_mN�Z��ߒ�ņ���N:�}V�3JM5wI�K��"��B��xE�妝�I����`@*6�7u%��ϐ�� #���LϮ��.���yI��yFR.2����3��阂��T���� �o��v��᫹���'���l�/f��_�Z��	�(�^{c��+F�s�@�K�ր�L�p�u%&�Y�eӇ�M�H�˷���Z�dK��K�e�?唵{&L2@��v���7����B%�'ř~3t"���WV��̝H6M���L�n�i:��mW�]Ŏ��f�����Ue�'s*qP,Zd
�w��ӿ>�Z����Mh.`�[���n��b�A+I�%�q�2�̖Oq�6�넝5��'�rb����v�j���"��Y۸f��s���z�t;[>n�������w��޾,�byΈ��a�{��)l�%~��l��|�C�������m�� h��&ޚ�i�1;�%�6�]���2�c��V����d+4��l����v���s�(q�V�rDQ-㼖�&��JC��}���|@X��\$��1}gհA�����?��/Y�6 �G��,�����_<>)ذ��cC�1�R�<�(㣔�)��ڨ���Tlj����3���7W۾���T����a�{^2yF3���ݸ��5�Ү��Wmqq``>M�����q�+(��FG��p'�ռ�͏>7��C<B�����oods:;B����/�k�n�`ǀ�k�g��<���31Ǣg�Y�X9�@�o~t�f���ғ�������T���Mx��cж��!�+�ֳm/���|��fP";�Om�W��������pLK�~iX�+�#q�32eY���@�H��d)��o�@��0��'�������*جxg*p�A���ׅKpȠ��ӻx���"��&��Oz�D��j� �=����t%��w����Mݑ�Jb��u�<�n4���"
G�K0�\�%#��W�OF��:_�>��>�D�2��aU���3lP Ǻ�hy ��$����Gɦ��|5s��,����=w
Q�"��C:�ZUNbAY�
nQ2���	�ѱ�q����� :�������n�.@;�b���F{r�^�x��A�*�l.��PB�Z����%���S�`j��b���n�W�$�p+��qpo��}9������Oi[2&�ns?~`[�����`b�W@�wP$|a�!�
�"�!���dkO̟�_�$:JZQ3�^�1��s q��£�(^��'Ctj�{�>�ˤ�:a�9��Ŝg�J�fs��5Ѥ�3=�����-�	��R������q���/"�nH}����'�;'��!yV�`;Z����R7.����f	���K>A�'^ +�S�,.4�+K���X��Ó����>tD?��I��Dm�6!O��w+��a0	]?Y�6!��+�M${��!�dA���n��י��>���՚i�A:���_V�Nn���A����U[�E|�t0Cϻ�p�b���\s8�+O�p��֩�7���m�J /��B<!F6yv�=/�Z|��n�B�Â��'!'�H��^C��o��i��O�9�uͬ�2�}y���2��C�	�F����pvF�b$�x�ns��39�K~!��볊���Teݬr\��z]a��EM������m�*�|��ޓ�i��a�3�(�;F��L�*�M"���)�jU�ʌڑPH�^S�w�P4�_�����|d�0�;}�"���|1�a��z��MT�)�cэlt��4N��h��t�R*�T~K�u)�7<�u/Q�^�#�Jf*�f>p�$rd��0`\aG�-�e���OԛP��^��&�zzI_�ŝ��@W��������Ǧn�B�(����{���h5ٙPǆ�U�K@zN϶H9�Jq@�O����u��]	~�����<��)��s�����BdU�=Ww�F[#�uҳ�8ř`�k9�q�āɍ�#y�KCRo&��9�kŝ�)�v��ƻj?���3�s�avt�AÏ�f��k(��N&c��D�:���V�O�[�q�{�'�v�V.K��R��z���T�#{=�S�0�zI�<1W�V��#�� q�2�M˻EtL���{��[CBn��J/��(ǹ#*j��Lq�W5.�|V5���ߏZ�F�N?�8B�t��>:�؏u�$�2d���M��h��Z�����L:�i���_��ʙA6�UYAϜө6Q�(4��wiY:+��.�'�=m�I�S���JD�����=���uW������^E��z=(����[�$�Rt�Q�U�Xi/F�?���RF	z��3������}��?��
<l~���k㓯ni����ԡ�CV鬾�jjG�?
=m16K}K�4�C�K02� ���4�1	�8��ƌ���݋�n��QU�˭*x� R�B��;���"�Z&����]�L�k@�U$��+�j��ﾦ�� ��ԞS�XU���fN-�L��쾥C�fw�E/�f:u����_��=�����aJ7�jh��<��͈B+x��f���#B��~�{3ӂ�s��µ� ��o� �1/��"����(��R��q"h��<N�yK��1[����jcG�kp`$L���AN��N�K7k>��N�B�1z�'�6T�s�1��}H}�}_g��Ƴ��ز=��΃=�[����ɦk����6�f��L���;��7d����lax]*4�Xk������(����T��d1ulN!� w��+�n�C���L�ePO�J��W�w �����@�n�w!�ƽ��_!IY�w��s����'EW���w������;��{�>P������Z�����3�5��VB�>��^*���7T�09i�ɠ�yҖ�?�|Pܘ������Iӫ���BQ���%��7����Id��Icס�|�JgA����3­\�𭟭����-R7��Y�p<'�{?�BKg�b!�h�N'Z�(R�l4|c�(����;�wY*���s,�ΰ����u��U��Hgh�6�U�����KgH�Cβ�S��2�^����׺� .��{RRO�"���
����I�8��ϵ(��X+q���P<a?�fĔ�Y��x5r9���<�D��ߔ�|���
�<?��L{$��PC�E��������^tl���g@M�	����t֊���&�(�A=�=�ˍ��l������!ă��0��;�$����%���0��5$�RK��׊ʘ�БA��%�
��!k��CM�ظ������!u�G�������c�sj��)��p���*{b���*���^l�S�T������f�R+b~Cdm;r��s��1(j5-^����1L��O�, �H��SF �Rn#I�U#Q����!訓aC'|!����jB��>]�X�r��Mh�&/1���~X!�5���xƊ��'���PX�>+���oF��B��ڥI)�;@�1#�ú�Qh�t����R�:������'Y�G�Ǆ_ڞ��'�:�al�a (����P2f$��(2Oʅ��4��lՊ���&+�-��<{d���m~�`�Ž*�<�ꇏ� ��Д�� ��އ��� �{�v��?�3�q񄷯��B�:�fkߐ���]�w��)�(p�h)���q#������=k/���!�G鲆I��_Q|���o��֣���YTu$����V��,�T���E��
�[�-��eR�,0Xh]鈻�n�q�q䩓�����l(O(^�)��8�I�&7�����Y�;��D[{@:�&gv��6�"��"� ��_�IV�Qa˽!c�rq0w4�-3r~6qֆ��R��5m7J�<G5fYO@vh��A��]Ϗ�x;�*�1}��!Sv�X����|�n����B�&dR�����	r3����~�`H�w�?���$��3�@1ɝ'�T<���n��a~"B���h	�tf�D�ю�� U]�^����2�{_����񦿾\eFǺ���)FMpO{P����|�V�ր�B�+��x{��Q�*�����ԉk����˻̺�ώ9}9Vj �xP�#��K�)�X��'HV%[w�a\\1�ج�N��G�ݧ��D��W���������f-	jz��l��Am&
�r�$p지�̅�	|��!0M��f����<�������%�wӛ�G:�ҷ�Yu�6�#�Ϲ�r��- a���@��O���N�i�*��gGM�`�5�6��Szv��P��E�N(����8'6A�w�O�]��c��Iü"<���L�=!���� e��ށUG�'ĥtM�k^<���"3}6!SՎ,I��C �%�&�!Q<�۾�CU����"QH'��Qy���e4�p�U�Rh�������W�	$k��5BY9J`���3O}7��q��	�x-�`&Ѱ{ӿ�8��6��=��9>�^��Ç�$%�<�Պ��F�9�n�� ��a��d�$6�/��ʙ�ە���'��,�Q�� �\�vb[wp��e%��;3���*�e0B�7���t��8��1����h:#9�:+��&i�c��b�I��)C�F"�u ɔ%��<��;Ο��hԟ�P��Z�h�Vq����˲H���,<Z�����q�hL��uD�u��-��p
�5!����T��;6(;�2�������]�'~
Bl�V+��_﬛[n�_�h��'c��:�Dra�'vj]�x�>�XċKx��@����<Xe�U�䣦,B�!CZ8��$U����.*�!Ģ���eaX_-�ۧ���������y�'�S���L~*��� ��]�yNF��Dڬ3w�w�J��/]�芤�N�k^:�#�����c��.�])M~�D�u{�J�\
�L�>�9
�|y���]5�e�)��K9H��D�Zk�>%(�c����~��jϒ8o�\/���ޱ�uµ�%�h����*�ae8^�9v%�.�A����^C����"F!b�H�7�9��P/N7�g���8��6ʘ���@� ��7�"�V_������E{@\��Bci��+�y��2e>H,p�e ,h��O�6>�!HTE@�����Bu"��ɘ�f���y4�'T/�����i(�^�뎊����fX�Md���)��.�e�~����7&��*�h4�et��|������9Vm� x����
 ,��,��a�>��5��f���Q1PndȉY|r�.�`��`�m�r���RR\gR!�:[o���@B%b{��dT�1Z�b��X�=�Hbֶ����乬O�������a�ԗ����P�@�_�@����h�>�(S��Hm����q�@�Q@>D�i}Sl^>�i��U�?Cy��Q����� G��F.B�"	�6�?*̓�
��vX�b�ܮ�P��݅»��|s���5��Â��u��<��{��Vs+t�;*MF�b�Bp�e�������z����(J9`�[�_�=����u���]�%��.	ə-C����St�������	�Z��x�����̖X�k.q2���W�s?џ�DO�!�l�1>�7���}�/��� j����N�=�~���4�A�t����+a�Bm(���A���E{O�,����g���R�r�;6e!���U� O��`"p�oL't1P̋d!�qW�|�pm�e���D-=w�ǯ=�N�Eli'%l^���J!k]���Q�Z��;��{�-e���I�~x�cS{���I�BJ�k�/�`��Z�
a�,qӹ_*���ŭ�Q���z�qr�>�:���ܷx�3�g"��$��"�~7\�w�I/u������Z(n�����,�.�-��}���̀w1eں�5,�2���X�����!�5��Jd��?	�--���w.}Q=6>�V��5p25�Zػ�"�{q�*t�{�1.@��а׌��������h��-�yGs�_,�����m�h_{�+�y8A�<�&*.����/;��&�+����Ly�!�r�����}n��Y�d�\���s��fp�j��Q�kB t�� �5�e��C��.5�'����%8���f=rݸA������Di��B�%�'�4XF��Ė NFsKAR�A����l/D�􄎒d����G�N`������� ~�����s�P���P����ĲQ�D)E��C�\D���C��)Y��eU܌�A��1֮q��|B\*1#-
Xi"�z�]a�9���/��B �4����R���Y_*8��%]�紀��\ں twǞQ��}�4p��F� �n�Z(P�I��=&��bs��Ϙ��.#�.:>M	_���@[�,H"���n�ey���+Í1	�%o�3m[���/2�Y!����=��V��ic�����VVkg\��2�,g�.��gd��1Hs��g����O2}�+X��Cj ��'/���0|�u���e�?s���C8P���= M���vx�&C�K�y��E��$��=R���ұ�ם�f7�&��"$I���pw��G�d��.�)��h�U3�i��u�l9_@,�����6j,�.}�r;�:늁��T}�7��0A�Ys_�54�y$co��nE�[�n��=~C�(pW�x/�R��!��4'3[������a�̒XqV.M)��Jud^�˷��M���.��?��&�����X���2\�\��S:9E!��H��a����[�SȊ�����Xp�� �%��D���m[���+�X����Q�]cS��]Y�� �)��-{�P��)���"�}�덒��@B��?�oE�VS��[؉�#3�^B�-Yۼ$6��^��q���������2���m��"!���7 DT�`:��m�(��|�n�N�u��_WՊ�b��^���;ѷ!��ڴIl+X���0��NKԩ�g^7�E"D4��<4�� &	��K��*v�y�f�P���fh�c�[����.��t;a#JDF)�����~��R$謐ߛ���6֞bugq{\D����R��T�������B�r5E��3��V*l>�[�/_d�'7�/B{��x�����_D�l� �hJ�Q�v#������P�����ZQA�߃	J���B����{~6o���m�[�lj�-x��Ά��:_R���~R�C�Ԍ�B-�/�"�G�N��s�W���ޓ[M��M[e�/�M�A��X��{j]���E����~[� ���2�UZ�^_�v	��\?>q�� E�t�֒�ܡoyݏ�k��T�f�MU�q��#�]
�]~����3�ϜL��D%��������k��9q�X��~�A]��o_+H��4
�T��LXV����V��T��L����y�z��ɨм$s'X��P̥��n(Ӳ��.�D��KV�ͫ@H�q��컏b��׵���*gݭ���./�]?F���EM&3��!����ׯA�znP�qƽ�_��6�t�ϊ�_���]�Y��H<�~ț/�v����b��x�J���9)GQ�8$���`�5��1@��S��1v��dj� ��%�%��8�..Q�>B�vT�����������G�������Ꙉ��v�yX����`B��N½)�9o�ގ��0>T�h�s�4^ǳ���A�0i^�/��]��G�{�G�1���k�K,)L�6�9I�u(쁭���~��M�k; ��G�F���֊��Y�TνaV.��B�UQkw/�W�KtU+fP��T8��ݣ���O��k�Bl�b���?-�j6���g����L�y�}YG�D"����zU'���s{]�����$5�9j׾����bDw��47G�,��B`��R�H{˗�
��il:7�+��q��@�O�	�ӏC�~���g����˟�z��i�2��wG(��h�'ã']��:�0WQ�Y�Jw��2o6�S�DW܈��̽0�A� �J��΀�uC��fy'��q ,b��.����U��B�0�P����� �xTGb�����o�Pf���=�(�
I��Ѳu��JBʤa6��W&�:�\s���5^�,��(Z���"��%܇�Uڛ�2�������w�����y�͆�co5FC����=֚�^~!�|Zl���<��.�ꄔ��� ����9�8��&>]wj�= ���G��Ou'����d����ّ"*�TC�O����jk<�d"-���8�o���@@t����D�E�R���zP'!qD�d%h�l�<��|������d!_�Vt��u��X��wlC���݈}m�.�<��/��`��Wb� �ڊ���qs�4���{�����U�܋QR���v�eE�/s���������li����@�9�)���"�H���������dL�u���(��y{$�Gt���yG%ъ���>��	j��yӐ���juB��`2��L� &���gkt���g�Ѓ;��z��ɞ~y�z(a���y,O�it4���N�o]���	�e��i��T0����p��G�-�L��;��(<!�r:gp���h׻�o�6&��v�0+1^��]L�G��������w��z 5^¸�̋�7�`��Ş"�T�b��������K[�	�S��D�a��n2z��5,�a���|�O������A�G�SSt�l�h�wq2#ƕ�Hx1�ldVI*/ԓ෭��S�3�-tĨ�㊖@�7�0��R�	��!���7�A���l�!�#�6�����^���[Ï>�aW@��)U(�_��e��63|~E��b�{1��=ӑ��<?+�;BR�
�<T��(9��:�Ă�
܆���&]#�C�n;
�{C�nDx�V�K�յ�d�~ũCM�c��!d��V=�h�N6W��ԋ2�Ke����^�E�u޵0P=}���츙�c\��CZ�m��U�����.0y�Po�!�5��ڐXf�� K|�ԃtM#����%[�e�Vj��5���5nDQ6�`4�;�i�r���֞s�T�˯�*!�B�[
t�ۚ*�iSB�Ԅ���p���5us�2��w��qe���AЉ��H3��,跥'%A}�Wl{��tΐ%��,�H]����9س�6r�h���@��_4���K@k��Ӿ�!������}[�L���5�� A]
SD��wB���q��+$�h�M�[E��W��^��..#�2�Z�'Dp�򊆬�dG�9�� n񮼈�"U��ۙ�^���m�͐�!R�Е�o�!;�cg��7���!Ӥ���m7;�!%#��� CL�T0�Q 6�}�7��µ+��e�3b	3�h�w��'��h�����\u9D��m��9��f��P��VbD5�J�⢆r0��ό�׻�G����$�+��0�i��	��N��M�1���_�xJ~��'3��zk���q&�s�A�[�G\�1Gi�@`m���a�+9��nYPkT�� TR��tΕ�֠Y�F9H^�7�y#8X�t��w�pD��ǜ�Ƃ4R���*(E���Tg�ݳc�S����Hq��C�~ﰒ�q�#*����HmS�+c;�6��Zw;�"�L��fނ�k�Y.T�R�|��L��8cGE��Pnz^>�)�ȕɰ{4�q�G�ꍊ�u?Dsތ��9z�dH�\���B ��U�����(2����=3�1:%��T��UN��K���{R'������}ٻ(��/�-�-AL�~'���cd�cѱy �TaȦ@��}�Iy�T� �P�\��j	�F,ef$�e�,�����oXR �ޗ"؟���L�����nG�� P�Rz�N��] ΀��q�I�i��[������"~M�T2$���3Qj3q\�u�{�;˃�}����_ o��1Av�_�/MQqR��g�#��ڈ{�N�R��z۲n���`�>�ZJ5�^��8+1����jz��fu_��Z�7�Q���?c������9h��Q}�z���c�poϽ��p�?g�6�;o{��#iԉ��j�V�p����������n4��3�.KW�+�a�w2it���nDfC��=.�
q�bPr5��;��������]��b��+���F���4��dP#�9�)���{䡆���7���/�(�Q���44���?MQ�G�GC�h<��u��KyD`�I���f=e�9��Z�e߿� d$��7 ���a�Җ��n���U��Qx<���\��3B�H;���s��c�z�h&�z��Z�8��t%js9�����r��H��w�`�j���t,ls�����X���!	Ě`������~�Q[�?H�������%dW�디����k�s������%ߊ�T%��k�3��q�û�U�)�O��GF���u����9��P2[��K��RP��+t�M�&u.׭٬��Yp�9ՌP����̀��4"�{Q5 t�Z�S�_��?�v!��dA�W(d��ā�C�Q]>�a�i�0�,�]s�<&Z�}xee�}���S�/Bڞ��[�v���w/'mvO���9��\���S�Pυ�s��-&��{���g|�b�R�ܨ�^�����g�m���RB���g���hA@��~�SiksV�=e���aS~ܾ�{hTsw���GJ<A �3j#!t"���פ'6*��˴��b@p�
`���@c����
Ԁ���}������+��'��%3.�۹��$J$�>�YԊ�o�D�`��5��+�@]���[/<�T�G�ϑVJ�1�uh���פ�k��57�g����F�K�{h��o���l^8#8a�=�EҜ1I]{u�f����&��*
�z��ȅ��wE�{���a��n�L�~7�._lbu�ʩ֥��V�1���{7S�f �:���W*�T'��7����%�MsJ�G�+!�.�&Z���]�3��8��-�%%�6 ���^X�$ٟ5幄t�p�%!QƋxv�Q���Jy[.]�Z�}Ms&�dV��0.&|B�t
�i�"LސG"R�z:�e��ԃ"\�dz!�����QMy�k��%"I�F7r�|���Y�)*��˵.��G���5������Q��9���T��q ��}/ar�#������N5ϑ�qa�Fk�0C9�j�2���]^�٢{&����v�)�eN�ut3�Fz��4���_�%��Ź�Q�:��N}\�{-�n:K����&����i~�Jb��a,ir��,2!px֠��E�1ԛAl!^b�����7Y2VE�5e�{ٴ��Ք$0�X
�Ӏ8��k�-
s�G�4�T<�6OE�sP�-�U�ʾe}od@q���	�@������B�˞:��4j��R1�Ē"��T�{�p�%�(�S~�`��<m-CE�S�_��R����`��+�~֔��6�bF�ߩ��������~��g��cå5qS��IM�E%�f����Z��{�(��പ^Q^U_��5"�l��idVC]���6���4w����j�
�SZloЄ�i�m�܌�:�=�:�g��˄,Ŕ��P�?u}�TL�A�r�$7&	?԰)oԉd���=$t
N��|.Ɔ���e�cf��&�q��qap�%ǂe}�9�1q�ܐ���X�f�HV�х�V��:�&�g�� �i�tO^>	q�)3��*?c�sЬ���(+�*�i�MfP�"D���A�H|�н�º?g�ԟ��Ҽ���6ҵ����Q�3��Ӟ���������`�4V��a���k��d��oH�Y�@w3�\��C[0t85ݩ��Г���Z$P���@Tp��0������6x�z����%_��4K�D�}�K��@l�u�{�2o��~W~y���G��l�|Pa�'�ȼ�Z���\���[�̫jh�G�0�����cO���sw�D��.ި���R��E�G�'~�{��i|��i���y9oo'��p��W��5�XJ��x�Fq��<
R��H�?B�8�D�����Φ�p��Ol�U���#��$ڣ"�(�m��O��'�k��|��5�!���e�}.���b�b�ZR���s 7�0��W	��-$Huۓfi��L}z���}�)Pi�ұi����������ERj���F9������p��oP����}�u4�%�(&�2Ӊ�'z0����ޟ�8K�	��a,!a%��]�����Xd���f�g+�ߖ8E�ѥ12o���%��s&�h��:CUz��إu�*ᛘMs�E�h�G!�<G�]Z	�
��,��Ĳ��vA��Ne�9�c��fi��?�Z�$���bu�/�)?	�,&��wBc	7FîE8���d�4����/��0�
��+^0tS���Ky���p��b]���/]Bk�Hne�p�X���?����	̳DnU# ��z�O3�5�$
T��Z��Y�����D��IC�F��P�h�_:���_��0�>�+b���`�^�]���-M������V1�X�Ά1�I�$g��XhS��a߫�	և(�z*��V).��K���å��M b A�����~FB`C�Jj�O�GMG�k�/��ƪ.zk���<���lV�{_����_��=��{\T,�������T��?C��ot-N�l�=�J�/��I��P��\DU)[-�7�a�Jn�{e��H���<TDb��[�+�)i�rt�w�pDO(,��('i0Wq�bQ?TѦ5��`ev���$m}�bvл�����x� ����P�m4wq�ז�܍mk��l)if�̹n�O+�e�\ye�+l�M����B�]I�Z�����-�ww8��nZ�i�ߒmay5&|	�o�bw��*��L	�&�k�]L�*\��.�v|��vy�+��7���b���*�`�T�m�P1KjQ� \]�/'����(|B�~�)�5����sDD��y��#%0�&��f�ΟRs'��l�YQ�P��b�#Ww[�uv��S����,=]#,zp�E�I��L�<����������w�k�3��vK@�V-�2����F��v/��J�zZ�\'w��t�5�Y�#����R�"��P[N��0�
KE#����n�=����@ ��1A'��!a�H�)}����U^ڎ�d���Z�Z�1W8�!�o�]��0�,�vR��F�Ա�_m_eǍ���6�b3�}�GGl�;�k�p��ݏ�(�
0)rr@r;���<�\��b�`Hg��[/O�8֛�T��5[���H�=)Y�P�H·�Z2��3�- Q3[JTNЩ9��%qcE�1���
�h�t8�߃�����(�(ӹ� 걩#�a����t����Ԓt�&��6[�KP�E�C�g�4/�N��b��1L��޿ ���{� a�9PS��ޜ���r��D���Dv�j'�z��a�6+p����醬`]��9��$��=+7S�����
�Ю�U�-WB�F�����[���ۻ��[n�E~�$��荓�ɉ�Z'P�nB���~�sC
7�&AgH_3�869�ؒ7\Vw�Z*;��z����e��� "R"�cK}'x�A
$�	(��[��ч�qn+	�x��3��R]U7�%5�����]��	���l*�.�[|�dr5��-ۣ�V�ğ��y�:�,�P�G�|f�C����p��)�w\�F�0"1��D�+�z�%�_�h)��S�ʌzkVQ���^nɜP����M0�՜�̘F��,ٯNȸ�{��6Q�0�/u��0��W�	&�O�e�
/۠r\�s�o�6�����~"p�!
���hbq�l��#��a�lE�����*��z�V��^�	�Y���ې�d�� ����"�B�Kx�>� ����������
b*Z&x����:�s�|��ܾkAy��Uy��9�`���ϕ��i�+FX���Դ&�����(,k�~z{���f���	���)FՎ]>��v��?2W���L�P[��N���B�t4?(��I�{�0�������Q�1.�A>��۰v�.���,�]��f&��-��H;���Ϙ�1��������n�U���˲jU��}�o�C�t�+�\�F�Ny(�_c���K�p����2��q�����̦�<P���	����u���y V��զ������G'�E�7=�e�G+q�1o&��8:NB������|k�`����:գ,��$Nu����Q��R�A�6H�;�~+B1�w���]�K����U�j��Ք�30$g�e2��E���%H����Z�:A,�×��� |��@�1�jۍ?B{z�.㱲��U+	=U��3C[�D&ǡ������2J��uޏ:2������&}\�-Hj7�wZ�DD�%����x`��%	T�֨,��۵(I�	�n����wK��9����{��������e��pZ!dh6kq��dPl&�<�/��вB��h��Xݸ�~ķ,t:�WP�4)�/7�qe#���1�%'�H��*�V�r��`�f�>*6v��H��!
�D�m-����1�NC�$�����or꾆j��!� /��4jcN��7���=�c�"+���r\ui��O`W��=��38�7m�5ԡ�ؓ��7Zq{Jb.���M��US�THNr;6�_�k��h�j��0�'VP�[k�U��4>"�<B5�B�:���@�0��֑�4��B*�d�Ft����kW���_��R��w���O��p,|@LO�A'��F�^,��O}w�f; ��7/b�{�5��BӉa��x!��QDP�i�@��f7"����pD�l+�m�<�vBP闇��r3�AN5�I��r�(NHK�b@�5�=�]�*�ʢI~����(���I�����| ���-�������_��1���=����l��W/�aH��G&m �����b�7n֞�V�s�����g�व ��B���l��JὌ�Z���D�]���k��gvg�t���K�D�#�%I~��բQw@(Cc�H�B���9w΃M��Dݛ����{O`����oz���v$�%�(�Ǣm9�b7��F�]D(���gR���BQpG���!y}�+;Z�*��2L����C��ɢ��^��)^V&]�Z�2ϨW"}�|^��e����O�I1���5=�Tg��Q$���4�i�q�ߊ�lr�<J��k�:�}�Sߔ��e����0w��T�R����� ��Z���[�T����Y!kK<�o���6Dc�&ڐ� �H�d%�w���� �>(��QH:-s ��_���Uw�����v8�d�A]���AZ8\��	���`9?Y0���x�QL�`b�^L�0TaDr�%���Vjn������"���JrSz?<dg�x�m�X��C?Su]G'��jN�}�ñ�)�~U>�G��]	9,
 �����_��5��>f��"k �Dŵ��&F��7	u}�d�=�2�
Z;���a(���
���R<�-��4�6��i�U��A�M&?��x��7m��P���E��+~�������pț|�%��?(>$|��ֹܺn�1_5K��L�����7r�AF1g	���c�+E�ߧ����7M�罈Xd0��+�W@7��T�o6RI�D́ S�'����%�P���ٹ����!�O�+��gq��,��n����@�@z������5NǤYqz�0�!w!���5�(ƅNHt����!G��woQި3 >����}��Zp�݊�ר��]��lZ]����8��N���#<͝���5���e������㡄KI�~�� 
�頂?��9��@D?� /[�/�f"S�}y&v9��(7<�a�+L��e�ܩ���$�����$^�y���C�(�?�����k5:�F %/���w0һ�'����}���'�s��W��|?�z�*��U��w�N!m�����ćf�"b�|�2o��� +�,��T�r:�Khͩ7p\�EVw;?�A+>G����1i��ۣ�]`��:7w��4�h|��	�m�H7��d�]�7|Z��T@Q�[d���~�L��Z*@�aas�c�F���H�f�=��-^��'x�Jy���S�ޖ�W�}�A�,SJ�_<z��1�LL�� R�B���Q�>�g��g�$2Y�.�=��ҵ+�;.�~�'�Ж_���
W�5,:0��z�y
|�;����c� ���8��?6��'���(m/�m�V9��:�vi�?{v�Y��#����+X#��A���,/��`�/����=2�B�e��*3.㒷ͳ�@��bV��	t ��7va�	ݯj�;?{ܽ�mҭ����hI���T8��BD��v��F�vő*�V�1�l6w��)�N��80�s�������!t,(g��s ���u��:��1BkC���{8H�^��[
F8%�7�`�G���(?�9B��.�􌯠��W�7,.d&X	t�R��&�ZTtX|�à�kl��|�}7�~�?Kj��y(���4`���W���Nf���&��;�Qb��\��s\.@��D�
��c ���G��;�0��)�e�q�B�w�I�K]�Q��ׅ�vJ�Q�&��f��G�r��T� �T��|r�������PTQ�^��A�\���p�"o�cK,ꨮ�G�Ẫ|�.�ߴ���`��i��ZP���� ���W���%8�1$?�&����W]gPP��~��m
r"��zn`&��z,����'o:�,C$�����'�9���ݟp���<57ƅ�
9͐(A�.���i�<� ���̝V��G(���_�hC�aϠ*�k���I�ǝ���_lr�V�E��>��*pY�I)U�ޡ7��ւy���I�7J�WIW*]��!���V0��ȹ�!@1����r������T��
�v��H�k:A�}��_����V3n�x/ =��L�W�&hG�ZHKH�EQ�������zh�k;��wR�A�9I2]8��u�a-����Y��.��8y�I��D&g<�B�=�cΓ������B��IIO�^MG�&�����b�	�w	��`F皷8��<�̹����Y=o�~:O�m���|:Gb�+�lO���Q]`6�lp,�Eo˞��QQ$C����.�
�^]�f�������`��3�0T�ƭ2ǜz�@�Z��c�K�&�~���=���IE�[��9 �����/��7:��Cvi@
n;�'��i�by/2y��x����d"!�{�r�1���n>$�|�����y�����kI��1�')�#l@d�M"S����vDD���^)��n>$2 ��ʎ���D���D��Ln�!��o��4����XXC��%Ά��^L+�J��_���c��eߩ�ʥ��(L��	�Hq���w;MRL�e���I���m����mk�}��9mE�]
��Z �	��1 1��39'��[f@ݏ�����R^�K�����Aqb���i���H
n��$�^��J�X  �!�4���;�������@;'�m�--��7n63�x��T���h�k����\ v���ʇ�W���z�����l�52��	GB�)�ⅽ�[���i�!hѴ8~��2���z�*�o����FL��!����CY�yi�k�2�hko#
��B�Lu�����^#��	��ލ�&�D�UÇ9녔�P�Ou���/TSRpel1�aƺ qG7���l<d^�J aᄫy���~3�2̅Sc?	��ـ���ႏ��Α�k� ��[mC����\*��;"O&rzFj��y��8j�@���|V�������и���x�jt�s�\��)ټ�WL_+���>k�r���2ܘ��%~��'�oLSPڒ"���-�;?-�K-�cW�IrU�^��`��p�({8�b�4���@OD�*���L+��/�c�_
����dE\.U| �d����
ͅ�/K�y��%dpL~^+s[����4$!,��x��b��N池G�04v��Ҥ5ص��*#X�ϩ���4��:|]�O[���Ü�l/���6��H�41�#��n.A�4à�˓�3!���<C"�����?�k�^�vS�G��ŏ\��:��i�����@���xs%t�r����'7l���17�cǸ���R�q�T2&��ɛxw7������tU�0���A����n�F6{�d���y�g&���<s4�<�W�4F��8=����Hd'��� �9ॽUE"�V���x�V�����&�hw��G7��y���]���z��}Oe�J �G��B 5�֖n�v�z�q��p��p��h뾶�� �4l��0��QL�]�u|�U� �Em.�{�%3���YM���T�쾓*[��?�����B�hv�^+}h$E*o�U����CWw���o�kn5v�~��,�Y����F���z����RC��k^������ʄY�Fm!�ٌE�ǐ�?^\�K+!<>�Ӟ�@�n�u��m��z��ܨd����(ghY�q6Z�Y}+6�����z�	w��jS4w<�IMK���\E���2ݯ�m�$�t�^���RG��V$�O+��U=$e�Iku��\6�g{=��+���ѱ��+|��r7�ҭG�����ڀ1Kq!�N�2ڣ�<��n�[�R��%��Y���V1,9�ȗ@ɲs{�B��)}����q�\_�#Q?��
.���q��^^v�8���P�� .!�� ߇��7}߷���z��-)彿諾��f�>��!H�&mf1Oⲵz�s��~oq7��p�?"�c�PdT�"�]�B)����\h��Nh[��:8��G	�Ҹ����� }n�X���܈�G�I⛡ѯ�w��M��Hsm�%"&*���LƗ.i��~���5��y� �F�<�X���"`$���W|�w�\��͈Q񲳻�M�5i�#\	���M���	ώ3vl.g���Ƽ�>���vgI�z�$��?x7p�@�H�����~�'��i٫}�4�<�9��7xyl��&������Q�w��|�38�����A`�A�M���D���Su�L��<��]���J^��TuS�Ǳ�����z����<���͋��Ft�H�����"�MZ��@��swc��D8{���k $�MO�;дJ1��꯯O��w9Q�-�P}fӅ��Q&�yT�Ǽ����j�T�l8��ȋ��Y�K��q����-�k�v�˘p�}����{�o񺨵��J�e�C�ͱ�69'%a�~\?!G{еI �(�U�]�.,fM����Ȣu+�Axx�]�	}��Vc���]X;�` � ����vf5aTv��2�������u�?���SkO��ҳSi"���K���Ƨ2ͤ&Bw�*Kh����5��Z˸|N���?�"�WLܤP!H#ć�Ԓ	�y����7Y���mUJt�^e�۞�$�V����s�F�{��F&>��R�kT � kT��i�Χ("�D���ʴz����Bz��l!�w6?�J�#7�fJ� 0�&?jq'�E��`]-�_{*+�t���֮c��`<B�r�~&��^\0e�W�W��r���E[��3qn��Z��T+p��n�\�g:�;�fs�?{�-^SWW#9�5�T���Hh�>5���a��w%�V5�����Z�j��W�%�S�������+	�Z�he�s��!= J�N=k�aF��GGxj��{�0�;��8ߒf��sv ����	�6��cN�^�s��Do��J�jɡ��#2�J!r�yߌ��X.o#�6����y%��x�C����i,+#'���a$�n��?�s&`�)�i�m�{��dZ��g%G�@q�����+m���W��]��9���:�27�*�s�
��el5L� ��E�f'1�\FQ9��PX���J�,�� t̐m��Sr݅$bO�d�g����A��(�k���H2��'�L��:�k̼��r�	/�R��G.b��r[�BP��ݲ|�ଲ����&l���F����l�'�%=��Vl�D?�l��Xt���t�h�Iz��q�V�>ǽt��}��ﴝ/��B*-��lPc��Aۡ���ީ��ts[�<8+ظ)]��`���K��X�U���0`Lf�3M�{ f��Bm��hq��|EV�Hn��AV�����Zbx����*4ԯswI����]�fU�Hw�	wj6|�Y�ɫ������"g2w�6���~L�]�Ҵ%�
.�p�w�"���d>�m*9^Pqb�E!^w�9Om��_'��H�Y�=���5S_#Y������A1 ���'I\�/.@�b�GyD?�&��r��M���|2��60�0N��E$�LC��l��.*�]��s��;�ʠ����Ei1c���0�U���Zl�g$^s��k3H��9KӐ�]�rd��j��:'�5���olX�v��3���o�`x���Ny���IT��H����0��f3Ž������o%AS�+�V��1	e�74|��W���`a�D�N�q��f�F�E�����GJ�:3����#O]�yu�O���NY��-�n�����ܷ�IqFn�&�.���wq~�,��m{{��2ǫ��H�`P[��2۰O�$㜁{��/��l�K�mk�]גuQ����������zl=�܂����i��� �E�\�m��rB������/�N-�a��������]�*���n�6�`a�r�+{w]��"��ڣ=�l��56��!�OB�g�L�8D~�I�Tph���H��qek0����[�8�\"���-BH��:�E-�`4�D1�塃�s�Z_�k%�y��G~����,��q�/j�?I�
��}V�[s۹*OY}ا�s�l�� pSo���f�OB�� 5:qSs��d���"�Z:��2�o�X�����ꣅjTp(����?�s��0��	0�0���Б�:%m"敜剛4f��>�.��?� ���n�GKS���ãj?cl5���!���������j���
�4,�L�y��Q'��ŚI�B\�oG���\��"���DHO������b����aE��(T	���;N+Nk�=S�m��r��3���8*ס��+vZ�W(f�f2kՏ��q�SN-2��=t=��j���S�r~B��?t��[�op(Q:-����(NC��ͱ�OO�U}t��5�����?�X��d�1y"�0�#eZ�,Ek��hg oo�X���;K��qA��ȅ�;�ޙ���?e�+:G|<#罞5��'�1������Bc�q�꺴���e�QNj��XF\!�+�f�!���5~>�4ܾ?�@C��G	J�G{�Ӑ���w���V���}�������Ƭ��T�r�/�K�^v%ːC���(YH˶�m���F�˳�#Jgۨ�c�f�x?�v�����Į�aNܴj~�Ȼ����S!w�AcJ���[O�U�q�y���=�Z�<��ڕջ��$�(�S����k9B7E"}�8�����b�"����3��p��BS5�!n9t5-n��[��N�rE�(35�.�Ẏ��C�dbl�?�������G�Q�{�������(���X�!�w�X5�����lOo4%��.P����k5@���ֶ�=�H���_R�$�?9�@�֪v��S;v���X��)�d A�:�b10���|��M��I+���Y�e;-��t��텰ʞ���%�0�&kf�8�c��P~�CiӎVr�D�^M ���G�o�?vN�5����o6�`��L{O$��)�5��=ZY���.`�[�9��ek�W�y:�j����O��0z2�-\)��v�k���h�ttY������䅾J�h�3�P����J���)�?��x��������s���I$I���B��5�sz�����I/ 
�zi��p��gk1�u���hz��[��/zOI���l�]q�1��@b�r~fZ��s$��]X�{u��� Rr�Y+�k�R�"�`r�!L7�����u�8�o4KW�rD ;!��iѩ�i�dBC�(����#I�e/��'��YH=R�좟z?6z(���S�ш	�u�'�Uv���}^:m���	����\>�* �Hݱ�#s�N[r����\Ԥ�%"�/�}冣��C{FR8Pf��5���/����b�_�T�
H5�/�o6ՙ��AI ?S�B=�od�.�i�׬"�p���^�'Z�s�YJ�k���bC+;���Qs=���9��%0�)@#yhBv��1ë%��0�����gUѷ���L1^=pԕH��|��?w9V�TN���(�2��OB<�$���1���yգU�I9w`S�鐬ABϖl�[W�{:FPt	�`�t��mF|pP|1���>��?c�rk��Pc_��E[l�/p��F���/^<�ܞ���bL��9��(Y��(�~�p�7S���T*�8��{��'D{����j�F�dr���P�f��f�.A�/�=<]Bȋ6I+x9���nD}�"ҥZ}���d��t�u�N����g!�Z���;��eϽ���{�0������B��R���ѩ��=f��ӭ�-Q�Bk��!0WJ�y I� )�Ǯ�+H��Ś�=��� Qxۏ�1R���[.��W\E�bAG��uȽ�<}�QjFmK*�[�O��4�"ie*���mJ���p��^��-2��ګ���ްv���sxN�~�XIG�ǂE�*��u�%�g
8��ީ?ئ�qOr� �>=/� {���ςp��nVز�����5���Ͻ�?�����A�(��w���h�(��0#햷����S�r�$}�/���e�G9���4�jF=�9Ԙ���Ifh�x�8����k�7�o�)�&�=h���s�ݷE�=#��*�3��i�JT�^�V�q`�UhL�_ganQ��@9�:�G%�̒��
�#������֬Y���lj�����,�20���4ւ$��y
ڲ���R�Ns�:*�0��
���)�J^�t3ƍPT,ﺉ�G��W�L��`�ZUS;a5P~\'�9LS�c���j?����K�����N�>�	�����V/������a�<.Hv,�(Qhw�L9�?�FE~����b�u��)�>l�ԁϣ�Dk>)[�Ͷ��/�c89x,�,?	�?D�����=U6#��Ⱦ�)P��Kl+���t���MmD**	���yT���&�(�֭Ek�{(n�%A�9F�m���(����`a�e��^$���Ȥ�G�*ܣx���1�G���e�V�ⱑȰ5��7�C�����L|Q�B��qs�[k�Phd6=��F�W�F1���wU8��n�Q�+��PWS,��v|ms�I��sb�Ͱ���Q_Ǐ�P ��[�U��xz�Yn�T���7��2����|���cv`a����4�ӭ�����Y��MR��%��ӴL�n��q{U�'^T��i�Q;����,���I�q�WR��܆<�>��S�|]Pt��NH&���~�{5���i�z�ZF�@fV}>�iִ_���O���@<hd��kT?�bԄۍ�Vf�)pp��mǤ�(vVz=,��{�>=A����n�	)�t�W�����V:>s	��+6̗�loJ��u2�$ɠ-�{R������:������^���O`<~�2"��&5J��vj���1ᎏfh��v1GU�hÈ~�Ue+�s휽��w�m�{ �f���U��0>i��"2��KԌ��]�ɆUk���^e���}k�*N��^ă�qCݘl�͎��f��\� �M��eƀ�TMN���U�(���~�v�bG_����LQ+�A\Q���0Ӱ�q�'M��sF@.��Gt4�����=�]�m�TŞ²l;F~�x�%YO�����\6�I���L�W[�Aֈ�P���K���"��?"��Zg�������uÔ���v���F���R�0���8�|�>�p���+F�WXK��?���f�CΨ��p��22ӷӦn��h-9~���#r�(F����V壬@X���S~-�J���q�B5�`W>J�5X�g�o����C��S���h���+Y��M���r
�}+�,��@9q�Ve�k��h�������n�G��=*�
O�5G@�fD�m��9m�ݷ���>�<Ě,��H+� ��}�V�cD� �����6dղ�O��r�࣮�Sw�zB���Vb�6���S��o���<s<�έD���"qԟ]0��#kڡ��%�R�IY@��&�h>�pl"/��6�<�[U��&^rj6h���@�#P�!���X��/�ĳv^�ܤ�Z3�	Ŏ��**�-�{y�K�F��E���;AyU�@q>��d<ͻFY��Gg��֔��%���]zk@�þ���R����v�� H�u�Q�U/8t�.-�wt�PO0&oZ���5��@�h*��Y;v7�jΝ�?R�a��Н����k%s��|`��A|w��!��Ueru��85�5[ �!��Wnטʔ�nf�\�E()߂��l��$��֕���P-�D�Wn�`�n� ���Fɹ����/$�P%�9Q~�7�p�Kp��V�?�@�2W`2Ϸ2�0�$��;]����&Q�y��G}~���f��\�,١l>!�W���_7M�r�E�����l�D&�&2�1�@�������`��T�/�#6Øɉ �x�`$��T���@�pr���u�2�A�	��t^4�y s�S|��`=oKa�w5��DO%=�Y�XA��Sì��9~��#Ȉ��Q�v�{�`'�N�%t�\ى��\>��������[�@"E���wO���0�c'�U���{"��"��q���_^�2n�垻�LSu�8S:�E��o��5��hԙg@��Z��/[����y<�M!B��Dd��J�:�Y\� h`
�,P�͉J��b(Z5��n�C�И-�)�|�\M�Y=�' F#R���*�8�����A	�î~*B�T牂ٯ�D�{�	�r�
���X�HyZ��T���[�-u�h3*�Ԑ��s�nQ����ϱ�Sp��5�~�yrI�72��?2'��~S�86�j��F�l�e'�ʈ8��h^��Bx�oۅ��8��@:�
�X��NS�F�f���v	��/��^��$!"�'s�+*�Б>O��ܡT����G Ycx+/�u�J\/�O����&F�[���0w�=�(Ok����Y,�7@��&ײ�_0Bv�*~����}���%��4|i.���)�a8��M*xOQ$?���ll�%X�l���|S�?����I3\���q� v�ĽK>�ܮ8�|܏��S���"���F�=f֬쳨��N��a`2,� J���j���J��Q�H1>T��b�N��D瘜N�wK!�g�F^�7�<l���ِQe�r*���_�e�?���nV���:K�ħ�����m���I�{��:`c��~�Q��%��,S$��Z,=�j�:����M��k�4�a����AO,M�C�b��ѯ���?��~4�x(��5�V��h��k-rBD�l�<4p���<�9tA�F��W�������
N뽱Di�ey��]P�%G�VizY�wO�uJ7!�*4*��%]���E���"�g������J�;�Go�otz�q�����t��Y2�u�:�_4'턍R���$'��Ҝ,��$U�13$m����͠#ѹn,�U :����:�H�q
a���*�-/��@_����rZ��!���(|�B��KE�!!�w��.��xY�Nr����);���y��#�)���������iB [���ۼބm�v� [�ƙɕ�ܠ����ڣ�G��a(�R�&00�r2�C�������$���Ɗ?�{�P�$���Lm/!�������<u���l�K\*,��j���@�*Sr��67m�0~���g� �E��]�ٴ��p~W
�-�6Φ�m�wY[2�����5a�m��w��؆���z�֏}�N#��U�"%Ym`�AR[�����I���#1���s�>,�Ew$�U����H��vi���̓��H�!�G��l����b���<x��ܯ�����T�f,T D�5x��#��������█D�uŰ֘��4"��Z4��v:r9
&��<�}d<�Z}ѪH߮է�>��D�S��)��`ydC� f���'(�>{O�"�GD�3Nj�K'1튱8�D�Fݓo�~n�"B�$���0�< �ŉg&�^ߐ!h�m����~�[X���:nzw��ZG�zus����dh��>L�#����!��t'���ϖoe%�P>~��.����X��6�wד�{�Z���Xu�Xd�
�X=t2�0���5����e����b%7&���0>���X��[�����D�Pl��E3Y�MvF]'��Iǡ2��O
"�Lh�B����H�ӿ��S78i�ƣ�;�y���[߱��<�] �A+��A�����U�0T�Z�Tśu�b��؈��6�*p�xse)��q;Y���b�[�z�T�
ƅ���¯�j�U6>+�sq|k~�(��z���Zƨ�w�r���^��>� c\�y���+L1w�P�g�N�QYN�&Uy��~'-v�P|���"L�;�6�m�^���}�?�w�fv�E/RH6�d� V��xD̲������U��B��o�n���>2�F(�6u� ��+X�)ɮ�|����/Q���֍��}� �J�s濺v#��Σ��ԟ��'�p��N@�3���c	�e=�J����w���E�`��������a.���穤Mb�G�/N�"UB��<��Ǒv5����K��& /�
�����<�F���Ww/v nb�7A�ԟ�KM}�83����b��k�⋀9J��>+^E3V]���{7yq��蹥6���p�aJ$�����Мu��-}]��yt�|F��D������9�큮3�9�E���d���T��W��fe,' �S��DdvATF��Wg|<l�b���(X6�L��{���L����h�4hm�V_Y6xTѺ;1�
���NN���?]��M!�ߩ�g��N�S&�LTB��p��>O�:������d���3�k��b���qIL�P6BH<��Y�q�������Ry�ᥐ���u�T��w����0У���e�h��>?q��KW�NA���J�$`�8b��4���Zb@�[��OJE�IΆ<�/�2��zpӲ:��1o�p��.!rHUX>��p�܀�f��'�c8.0ְ�F|BԠ���S3A���bԊ��quH.w�s3T�/S�S�6�mO���I�C�ݹ�����O0�s�Vy[_D�͇�}D]׸t�C���w-��r��!Cy���y��z/4{n�D'�qt�xy�x�N
6�X�r9�1�w�!/���у�JOh�E53�o�i�SgJp��/;.���;#�!G5�ծ��(�۔q����~����a����������ށ���C�ߋ]HM��b҈������1�o/ޜ`�X��
��3�g�+������I�@.�>zJ�*�8U�,��ߠ�K���z�c�p�ӡ���Һmh��0�'T���$B��ԘS�*oo�X�z�@o3��5�0#�ҩ}�?!k��R��@ͻT���zZ
b��Dp�{�<6VD�5jЋ�|� ���o4[:����1�t�@$��C+sڞ:���l�G�jj�y-�)ӊ����4�@69�Z{�Zx2����,/ԘC��"�q��1���'G�	��o>��DQ75!����+r�0V&?��A���ˍ�3?]�	���}���:�E�)Ě���XIۭ��i�"a�<Fׁt��'�5�O1����Ӯ����\"��#R����ָ�d1��+���@a�eG������P?$��p)��^P�Ϫ��8��ٍ:�_=���6�PE�����k�P���/��Qc����2t��o��c~�D���7�U���|�oUY��`����;3um���aQ���@ڶ�<i�x�t�
�`�$�E�(H�(�ѥ�!���_�+RH��%��$�yt��o�H��b2	6�����?EB�&|Ӧ�3��8h�KVC��DE� tQP@�b�C�ڰO��w�����g�{���8�G�G󬅶k��	
���]\2_ޥg���/݇6�����`[_��̢��*?PyY�Q��bp�L�Z}"k�p��ީp��Ӧ�19�teF;��}%�k�ޓD�d�� �U(��s�+��KZ������'�3|��s,`���6~�8�?l=<
�	��<����H\٠)�a���� 
�K)��/��Y�����
Z3$�$��������T|X��4V�yg�#��k�C��xW.�7۝O�"T^ 8��+�B�^r����ƪ���@�*���a���Q�u��n誙���[
�O3����-�J-�g�T����Jsa�D�ኤ*k��\�����fK�*�����-'��	���Ө���r�W�v�,��8Y%I� g���Q��1-�Ɗ�k�O�"x^9ɂ���\�38�����V��J�Mu�流.�|��GL���${�pJ��ɢ��;��@K-�����x�9��.;J��ꆃ~k==�Yy}<�슽�~^��_w>���]���5�M3��p�&���Bw>o�jN�\SB���׃.�P��G0��v�nJ)��
�
D|��˫l؈\�l�ߥ?}��K^�{������˃V8�����|��gRq��dߔ9!�9�{*�������	J_8ׄ$�f�(c����&vT�+'�@��8�1�q2GO�+S'ec<������k�ycw��o�`Ԯz��*^��!��V�Lj.Pgr��p������������︔�
3��)10<�����AN�Z���r��>
���-@�I��B~ryK����$Z7U��������|�Y�z�����^�tt�����D��5����n���$�w%����K�rsA"vC��*�C~ ,Fz�I2������q	�ej��iA��DD�^�q��}�Qט�-��e�[g��w�(�7��V��J�gڕ*���Բ��Ҳ�]�V�J�ma(�����ؙo#�,�Nt?
�=:6L�@�#���\�{��q�:7LSwD�0v	�ɼ���},�}�},1�R��>��5>V��>�"60���))�Q.1x�|nA 7�ǻ$	D�~���tl�T�L?nd�,E�¡v�wX"�Ji���[4Y����d?4/.��H�ΥdU➚�閨���87�?%ׇ,��T�GV��O�˝�7��C�Zy��)]g���/�H��&8-($����Wza^ء�qL�+��/ښ�?8�D�劎�8��#��bl�=�(u�`�Ô$���\モ�x���b�X��4�v�lVA��6�X��� hc, ���4W	�`T�֊�2d4"N�����2����4���%�5�
K���[����hG�N�k���'�U��� J���'F�D��ZK����i{;{���a�Z

��Fz��4���ܣ�e�9V�	����$��VÀ�I܄�����B����ԬΆ}n}"�|�z/gڴ��hE�� H�����F� ��|	�|��hIXE���8�ӳ�+H����\��&��,>d}�(��"��=��#�X�x��;*)k�P/fX(�Cb���U䷖/��3��nZ��l*d�#h(�_�K�0 G}GA���]���	A7[�}&������I��dMu�{V�+�3�z�C��yDԦo)��}����[S�H�z`���"U�bӁ����(u�3���g�X���P��������I �y����/�s�^�V,�Ƙ{�E��0�n�<�����V�]�|��``�T�%���!��k�
���B'`9w�W@�4w�vW�"ɣ��:㹼�tz~Qd���H;����kI�m`sp�e<U�e��w��/b��G�Qꝏc\�B�`�Bw���.��hN�ĩ�c�I�_��BTB�ϛ�j��
����S���|������x�?B<�<8���ܨ�*׷vC#ixS[o��Z���l��x��rT�����V6d�$��#�������h���C(���Y��86κsQu�M�F�Q�o���c���xjh�s��&�Q\�$��lO���q��P�K�"��8��n��[TV,gZ�^��
m�5��L%*��%PZ1\ow�d-����nD���1�zlR����8���핉Z���ŧ5�x��Œ�h,�|�UB�mp(b�+��g�����DwD��.��mq.6�T��ltX5����F���G$O-��YwR����X
�b���x��'���c�-��j"��fk��$mT�S�u1�͕Qmn�X��1�b�Z3U>usD����.�8��j��W�ȹ�O�������e�%[wsl^&F��Q�HP��]��Z6ɺ0q94 ��\>�:�,l��8�A?�m�SU����G�]�&�C��,����c7�4�jt�� �_��xiI��-߁%�����"���#['��O���*1\w��B^5�A�KV����I�åVZN�ԒB�ߒ��X︀�%��?�@����j��M�2�*�>l�6vs~���J3pZ��O�1.�*�P��7s_!a�8�2}���S���+˗��)��(���˾l�6q�K�T�(q��X�L�x��ޔ����c� 7�O�hɚ�jX�D��|�I��\�Mu���8�Ζ�{�^9��LK��8��!X�G���[�<���HVx@\�y���@����o�DOM�
H�$� ��Tåf�:;�֭;�K�z���	�;Eޛ�d��:�Q�����6�-Ow�q���f�@r�ՊL���	�,׉�#l�Z$G����*-�;�P���/a�C��v���M��\�4o�)c��5������d�p�OTgv��hZ���+c�78.vs�����{m��U�o9�a��ZU�i�~�X-݌��
��l#Q�CMTC8�R<�%Y�K�l!�v	�-�J���"4�;��&^/���d�g���������v��7����>�$aj�K����"�B�/��'y72��� l���
��`4�sԬ+r���v�#�>�
��W�5@�����X����K_B�ѱ�W�wƚ�צh��(!:)��>3�\����I��q^2#���5]OFf��}c��-����M*7~�����=�G�����#��e�C7!���2-s���U����}k��l�q|�S>"�4Q��j��6-�Ea!�eE]���Y�l�:�����9&8�b�v��ҳ�Omau8��4[Ϛ�x�T�O����Ɖo�Cf�m]L���r��Z^c���������[t�ڻ���$���R�>3����+ ��.&���b���H>�;j��V�����ۭpLsQ�"�2�4��^�C.I? h+�պ7r@�/H���24`��_��JnF!r`x}��y�6�y����Ӏ�5Y7C�w!uѐ)���Z��*U���Bµ4���(�N���^?U1E�i1�&Q�g�7:~�XO[�,���xm�d8f IaO�x]X����i�7o��A�O�i��WÖ���:��{��/!0�uJ9|���e���)��d�>�[���\i)/�ݩ��@�g�E�ץc���s��Q�I��3�DL^��L?P�]t��P5��>��̢�P�Y�*�쳀j��t�B��!W�V�,w��@h.J�����	k�X�Dl�e?����J«�y�W��:�����D
"q��^T�Zś��a&��?ϥ��$���i���뮾i���M���F_thl,�Kp�ߣ�*�j~ӝ�?��*ca��m��=�ݴ~�`,�R�ʐ�J�(l1������kϹ�i�5"9׺Ē`;J�j�3t�¸�irV/�u�2�� �4Ed�ڣ�t���\S��c�'h�x=�՘\.n~�'>&���g2�ޔ��D�5s�0��˳���5ڃ�^ �����LHc?f�p����z�-�#q-χ=�8�Syq���qR1X^��z7�u�oe�?hƹ��+�3i^�.��á���ذ�O)Ͼ��>�,Yyy�P��).��)������C�&���C�{/��o����e��*�dR��6u;e��0������Cl��(��^���@`q+�F�@a�ĩX����V�Z�T�ͪ쩃9���m�r���>�G�U�C�x�܌�w�Oa��W{�Q+�Y���7�@&�df����E��Q8�޿p��1����s�|���� x��q�>�"%.ܥw�A4 �k��]7�9O�H���^����)�Z����ܺ�/�_�|e,�$�{�'l@����'Mn�z�E*��M3YFe�0*���r�_�G�םrP��H0C��������e""�����=g+\T��|d�G˷i�F'��v��e?G͂BLY��Y��J�a�)��-E�f_�jQ鰟ōi�̤��B�7>v  ~՘P�X� M;p������@��:�<��t�ۼ���X�%yt!�Jv�q�ս�f��>���ޗ`Q����r�E��>0�Xf�l��Jd��7H3�	�T�n�#NO'����.���?}���� ����49dƁ� �ͼ?Y� �B^4�<w7pV|;	Bh'LGE�wt>?3J���+)[إ:(%����&"�;N�
�6��[��9胝G�HM�b���.T��R.�6�Ӳ#����<��H�ȟo��*\����ח�z,]��&&j$��}��؝���}��4gXz?'x}(ڵ���'��C�
uA.J�~"0��m�H�:�N��Dd_�=>��1m/ԀlX��])J0�����}���ڇ^�BAb�;�� �c��[�U���>�4�$X�z����?�ł�2m�̅��Cм���N�}`�����o�ol�au�Z��p�(@sSJI�+I�i�a����!k�=�h�
�h�-��`̑<��h�K���1��x�V�e�c�T_�*��XG6ZlP�{��F���\`�R�E�e��A)�����T��5ýV��8�W���TBTx�q2g�i�H�~2E�!�c�*�9�i#EI#b"�#$jS�s1�c��d)7-��-�.��<FDR$9k�%����s;5D�:�(
�ō[���X��sĺ�|�Ue�'�^�cE^2r��}���t����)�����km&nԟVϝ@���i#|}�M���f;B�=��4���!O�kEa� ����_�p菕��!
���*�eox���S���KV(9�g�m��ߌ4e�!d�'1{�S��_s�L�B<1v�<P*P������gdDwq��^֖/w�3OPY�<w���D��G(c��" +�KbqPK�����W�S��M� �T���L������B<���;bu'z/��Ȇ�N����9�8mpGe�6Ư_|�k4r�y�m�M�D�������8CS7RS�*����Wi��ǋ#�ˠ��`//��K��pa���Y����d��!�{�����yR.�R���uP����9w��x,>��쭜g�)W��e��|I	�iQ?����h+�]�Q�ć����-���e�����dQ�*(���U��;%TH]���[�l'5+^^��c�/-������N�H@u�q���5�t#FU8RP��DF�4���Y=����:��6ߣ4�@�F� ���6��r�p<'�|�UK�@�r;x.�NWp3`�ׂ��|��	Kˁ����ma�Qٴ\��q�!�.����\����{�2�e�:���@�$���S>��>p�ѳ䱴k�/rL	��St\�����$����:�s&��ty��` �o;Naj���@�H�s��ꭸ��}�M��D��S_��$}۷*��sw9��!����ϐ8�{�zOR؄�lP�a��:^GǾ��Rd�����,��%�U���sEt��C��Q����xz"H1�;���O����OVxz���xG�{n��(+'��Jˉ��w���b����P<;\� ~�Jj�^DT0�^o�"m�/���!"DU�:�A�R�I
߫���[�.�S1'��$�-��5H>tQ4�xa���|w��O����P(��$����ٰ�,W|6��֓ZL���3S�%�d�FZ:�"��T�H�,,��ݔ|��BV"V�M����Or���$pO�4le����O�SLp��i���uo)n�s�,MTS���S���#�43�ٵ�!�?�~�ƻa.���B�̊`�� ����e=V��[����gӤ��鑛�Jh�C_]�}#�l(s3F�b��!�ӌ, �g�!�y�n��A�6��^�U����jy�{K���J������6-4��*Z8fxسi��r�i�ñ7%��1P��&~l�\���%��O%n��zj@j~j󡊞����}f���C��-A�r[[���"�,XV#��C��5!I������������+��qT}6G�b�_��׊��)�ȶ��n�J��X��K����0��"a�ꪱ�@$j��u�`W��@��&sv��t~;�&ߗR&���}�0Cl��v�+?]ẃ����7=%8�����5f�x������E�v[2����ʔ^rq��+M΍$xk���s��M�Ϡ�60���Y!�l���#��}\��/�O�I}�aE�'�p��]�$FP֥!�5�(0n��|ȞEi��]@/�0�)V�7i�>t=�4��OgE�ŉ���K�P���(���'I*�J���(VP9�9u��<iar��E҅V`I��� '�dF����PNCq@O�,��3�N}�le/_���95z�{�LٶF����NSo�����h�4���GɲC�ֺ23H��Cn1�,ri�緃�Heo�'i������fr��u���%W�V*�[��"h��g��U]?�y�,�4u��_�3�xдSJ��^�d�J:�p�Ƚ��F~�>��u��t�{&�]W���"OW�*�!c���SZQf���kآ]�b�`1P����/� �Z4��QOy ݞ�ĕ��:*݄��v�s*ɂ��uɀV�=P�V�ڣ��Ѽ7yő�E5&Z�a���?�n�+{6��(���(���#P/����??�4G��(#�e�ӦaH~h�ݳ��5znq0�[��^~7�S>.eѡ�#��떘�t��ŀ,T09�Ӡi�z�8Z��8bY����UѯnIq��!������+�W��L�|n��Cz~�M��Z|E���s����J2�жfkC�ǆRF�V���~%K'��;p�z�y�/��ZY�ۋq��k���80�҉�YISK�m���?�?�����p�kbS<.�и�C�"A��Zk�ӦBb���!��` �n�Γn��$�Q�t�9�$eD�����e�=:~	h��
ЀT9!C���:L���ΗX�:�j,ĶQ�'�����5߉�8��<�V�(�y1S	�VÓ�clάN��ث��q>��/C{��QO�����@��9Ԁ�1�n��꣒��=$z����k��6��H$`7�roЂl�O�#l��/`㍯rD>u��ۇ��(�ǱͱZ6q�(���|�J��� o�j�wI�3�#��Pm�,�,<|X�v�6-��~ڬ��/n(�{d�ޖ�˳K�x���`�Y��Ɯ���c��-�.{)��`����i�׏͸��9���uK��u~������Cvs�C+Za�g�2ܟ��}�?��=ک�u��v/�����x���b+3<PR�������%�t,�b�NX�{�P�����`�9@�q��ŵ	���6d�����mj@�OPC����6j����?�i8���	׫G��guɂy�:1��W e��ƹFq�V�{�����n���'.MR�D���Tw�M�09ҽ���G�	C�e�%e5�.�/��z��j��)��#L����V�|��z^�����v+���C(kWl��^���I�%�\��t�#�(m��h�����׶��v�vX�+͚��B��	��?��k(Wb�f/:ш;�ˬ<�"l���P/@��rô�-a?��>��\]�`፩��'^����;/��%G%�'��P����4�؀d�JL�𠳠�vv�鉜�2�.x<CVpE��J�0f5�pi�ݭ�%�q�����R��Mͽ�Z;��;����n�H���dE�%�h#2h��G�순2�2�է�k+seP�9����f]*��]���LD�j�����ޖ��C$��v���D�&�WV��}#Gũ����D�]K�}��Ⱦ6y��;����"��%��ThZQvE�_�
��t������d���'U��B2��?��V9��1��R��Hb��kF{�뼗�I�^��2�C-�|�3�m�z����W�����L�t7$��q��)AF���r�gʏ&ńf���S�4p|SF����(�e�˷�2���߼a�����nF�B�%B+TiDG��olۘ��e+�=:wu�4#�:�]v0����Y�@H�D��>Y�E+����Ȧ�E�~�v��~H5jJ�W/wG2��o�`3��[%�o���_�
	��Ca�8BmyMPo�����%����\�F�Y wdO��ID}�*�Q'
aV<g*?�?�����b\n���D[x�%�"�ׁ+��.�"�O��uΎ ����tXl-JK���"F|�Ta%\��4EwP�,���!o��MP�����rbO�#�b�)���ٰU�:ŵR�;h<�,T�K򅓢Qɽ�t���?R]ؚVߠ����FU1���ڑY�-�C�_�*�ː��, �%M�g�)�Un���Vr�=�a�i�'��voPY����	+úh�YP�@Fݧ�d��a��\͓+3�7����w	U#�)<��I}]�P�Z�D����O���֦Y��`x��}��V��hU�A��LZ�s�qL�=�p���R���ʨv9&�bU�Ѭn���� ��xĤ��1�1 �>T'�'F���G�� {��� �^9X��y�Wj~��_�X���V�d��ÀPf�pRb�OZ	H>���9�d	�����(�d����`��e�h���L�o� ;�?i�����dO^I_�qR�A�P8�M<;��a��&e��ɀ�%yM���o.�A4��I�<�dH�YߴG���39ە�W$��5x�<η^�3�<�4���=�B��Ot5�̰�q��@�'�0uPϛœ���� !<��ym��c{���W�"���Q� |di/L���Yӿ��`��@�%bkͬZ�xP`N@ꩅ��ݳ�t������)OR��Ͳ��pm����A�{KpP6�pRJ|g�٪�g>�fjgK�x4�yS����O��)Un����%W67�������):	���>�h�[�`l�9#ü�?Ꙓ��jEL,xq[��g���r�Q�����ED�|?�>�t9r���B��d{����\��MA��Q����60�������Z~P�(w��*Dd���[�<-��G_��VLSGs�g�Ť��e��
���2��]㓾Jw��x��Ȭؘ��e�Ŝ��EI��XeFTr>���C�le��ս�l�YY�A���Z^�uZ�1+��Šp����.�i^�y�O[�]�aX�)��z�`]����P=	�$�b샒��\l����k��PU�Ծ�"f��y�طٗ�����b��6�A)�:�#�U��\t� η��{�7��c�v ��=��DJ&�s9$Q��Z����ȧ�j=�X��ޞe'J��휡7��}� {�=�x@��	������Ԑp#��|?vC�3�@rm�1����ժ=ԯ��qX�K1bW�]Ǭp��X��e��q��G�N�Vz	="?͇��;��.-�}���_OʳE.�Ntx��]j�A�f�M�l�	�H�snF�ה2��K�����������81�*z�#R1�!`�Hˡ�}���4N� AK������Qx�2��?�ü(�X/"��j't�6�̪�X�I���ү��پ�F<�j����"
���C������L��Gk47�f�D��g��}#�}�G��UŽ��i���)	we�"\�AuI,AI"@��ʷs�)��+2�D�^ނ�C^e�R#i�3��@�a?���{�	,�m_�>t����p��s�Ts��a&�	���ɐ�$����`��t��d�jÆ�|#�`M�|�m�n"<�!��)�Lw ^e�UE�%�2 S�d�6s�����?��h���R���F^�dl;(�u��	P�*U��>A��������,�ߺ(�Y"%���E��(rL<u�	��D� ��x[Pܔ��DۇN��7X�^��32'����	�&�����*�Nѓ��[�1�>I~���9�����R�@2�l��� K`V2
����N�>G��^�	��$m1�a>��5��7��,V7]<�5�x~~A�qw#��V(����3X�������$g�k��[�No����X��Z4L�+W��{_eQ����u�t�&��SP`X^��CϽp�w�: Qs�I�#�v\�M��0�ȫ�emc�J��iWZN�#zFd����sw5i�;@�Yf��Ҳ�b��00�k[�� �!$�@����j	[ �YAw+i��PE�b����e/�Z��L	�j�}i�*��+{��xɊk�b�>���,ó�N��wk=5t���N+xm0��s����0�`�1�;"P%�\N	���*a���a�@ਈ����߶���w�?p*ק����Ӆ(���g��Pnn�)`�0*~a��M_~TG����W,g:U5�=���z�7q��M��W'�3�Ս@��N3�y�w)^?�x�����?�>F�q5�o��p)��gA9��Y�e����y�0r��1��k����(�9t#+�I�&{��jn��DoA:KҬ�L��ʌcڏv�������鑯�E��e��)�m���S$�[�ׄ���>Ջ�dĦ�,�&�v��F�^M��7�I$|����E��s=J������V��
���l��X�U3~�,[�*uƢ�Y�Ԑ%b��8�ڻHh[!�)a�2^�>i��Fi�t��&��-{��ĤJ��Zɞ7�nawa���Y\��OX×{l��83z:v8��-��ti�t`DzU��K��<��y�@v�u|\����G
H��_Q�YZ?�ܑ9>3�R
�$?��P����(+�[PǷ/�q�5sŘc�
�p^�5�
��pH�}fO����6Lµ���������Z��Pi��2s��|�[�����q�7,�J7Xj�F���ŷ�K�AW�L	|��$zd��/�0=�-R,36�
�Ts���ȧhZ�4,����	�t�T`��[~u8�0#��>i(����jy�R)ۉc�3o���7�C�蘷�$�#��ʲ��w*ɅR�|���\1L�"�&�>k/�h�[�NuXnA7��1�3�^���o[mB�iIt��.��-�y�i�U	X�T�&C��ʷ�1Gg�܉5��%��1��������`�#�!�ۇa��/c�7?$��)���1;��8`���gW���왁�:�	���Om2u�g���0�`�T�X�"��YAb��/����`��h���,s�=�`RA��]�+j2��ܠL�;G��%-�#ȪH�3ћ3!��.�a�wǞ]�5�*��������o.�p<�͘Z���MĮ%_4|��UJ:�DQ��A�9�,z��ED�0��.1�Z?We�,�u���?v-��x���t���L� �1�f�X�kz��<ߢs�N�3�w8��*�Kq�r�g��t\��75�a [�K� ��ޜ ��#暼��>G����?�B��[�{�l��7|�ԑǲ淵W�݋�8�ke��z�F�ۃ��,Q~�A,��P5��2Xa������� �9�(-	�5������|M��y��c~!��]!=�X"G���ő��R;_��(3���0�7���瘙�-�u�:j��n j���S]�'�⨢BO����ZE�ݝ����/�o�R��[}�Γ,Q���`-�m���TJ��G4LY<% t�'���Vr��F�m�7���3z0c��,.uX��ᲹB��$C�E�O�k��T]��0{ȑ�%ɣ��&�'���!w���c-& ����t|<�c$����(��ψ�3$@H��Tj׷̝�dC}�ߏ*y�0rF�C�f#��_������u�W��G���I;���\���:�Ww�4a��)����a���\�˅o��!6�Z>�`/D)y����):w4��/�{r��u�ڇ�;��`C>?��I�k��eD�q���$��A,�G�Xl���լk���(S��19���G��^�N^H'�/�3k�s�p��5Gva���
�h�)t�ټ�w��A�W��^�ے�-4p��܋Y62���.�L�)��;�`$E�u2��Eͺ+Nz!��?�������<��X�&:�0厜OX]uJѮ~�=����W��oPrW䚷�^����pK�ơMQ��s��Ő�����s�I��l��d��fD<��ĺ��C��D���^�KT�='a^/L˦��C�vX9�L����:=���˘�y�*�%�\��R6�������Jf`�0��J�!�w �1a��0��k�b색	b\��5�7Vt*>K�=��5�����:K)�����*b���S�������qVu�t*�#l�g��>&�5B(IO�:�$�{-^q[���i��,d/����V��/�Nw�K�u�n)��0�A����l~Ct��C�t�Ծ{-I��}�q�U!��a���|%F��������c�a�R4�z��Ff?�U�
o�|z�Ӭj�dS�N��&�5���*Mw��d��(��{�4����ho�%%xf�ʪ��V�7?/T���N�c��s-\��z�N�`�N���PK�u�*���Ek&~��?.�(�8Tь���g�[��1I����.����
9܊�E[�^?K�8��m`�7�����k�z� �yJ�i����[�k$d�9��d�?;�nyx�hx��S�U���4q�����8��ISss�7�d:d�_���QnU���a�Z�JY,]��6��0� ��EB���oZ��j[}�g���<yV+�ngϻ|"���Yd/��o�Bא푥��.�l��.��v3G~��ԼSD\�.<#fh���u�Y��Md;�ͱSqJ��2��0F���(�dZ�z佣�G�v

@H[�Ti���h���<R�3Z��ˑ��ļ9bd��5���ula�<��s���ALV�Y�[0�W��s|.���\[����]�� �CqK̻��W.]�w�-vJ�*x�HJ)M��$0K%i�M�a"�8�*��E�xRzr�\P-�$����~����%���*�2e�����zT�R�щ�o��s��i��ʸ���Π�WA����"�'��fD���p)���s���L��.	��r��I,�V� �Ƞ��K|Z��� ��t�ڊ�기�\�|<Ӱ�w�u��$D���D���:3�܆���˴q��g�y��(�������P7d�i׉�e��ٍ���!UbtkI�Ȕ���*T��|wͺ�E&3|�?������O�z���K�v�OϚ�sqs��5�b�??vO��A$ˆ�F<�5�+'3����$�E��GVj��k�3��lV�OUg�n���ҝ*��P��X�����АLS���*s�oۚ'�$h��y�e'�=���EjX�i�cV:r�3�`B�#lmz��'����->��v�4at��yN��ߜ�B�����ܢ&�L���s>�t����'��:���-�_Ħ�|�C6cO̶�#D��� �#�f��_w�>UWEG�la�\#�4� ���M"�xo��m�+��U�l���O�ސ�4��Aw%=��_�fy�)��H�SO���7;)�*���6�k�����n�zc�S�C�h2emg`e���0R"�h�vh�FmD�!�`�97U�r����W�&5��bZ_3x.�(��ɐ�n�����|��;�w�#L���:�o���4G��;�C��M(qJ���ѐ�nz� 壃�3eG�jd�[��?/#(d �s�i7=8���D �������M�Q�?�_��s��L�K�f">��}�6k�a�i��n��;�M�b5��
!c3Ɋ�	k��+��ˁ��3$]
�F����6����)�9�!b0t]�s���d�&1j*�������&��r��������K5�N������˖�kr�^�?�tp��]���Y�J�� �� ���"f�Pi��f��A�7�׍Ns�l� b�3l���:k��]�V����v\�>;L�#pN.rxE*8c���z(�S��2�idl�?c��BTζ�]j+/C���܄*1G�� �ek� !�v�R��F�A���aJ�x=�<k�o&�����Bi�l���Ή�&BX�3�A6�C ���ş�������!PM9�6�)�����šZ8X�ߣ$��P�}xc�O�G|��<;{HsW����\<�`<�B
i�L���@�~��#Wd Nٷ(�0-m��AB��.h�����Df��V\nq�)A�8� �"�%��DlV�˺)�f[6>�ϣ����B�W�E�\��:�'�,����\��?,$���8D��~�
i�	�4�.�u�ZYN�~G�C��'1�F=ְC�>�Q�z�mZ(Ȩ�(Ul�v�u�+�c�Յ���MߞB���,p5��QF�f���m����N����p����笰,u9֗)G����bY ��ClyS��Ճ��6�����UT�Y Q�r�5����;��X�< ���LC���kZ 㤓>��8�&'h�04�ܗ���K���ޣ����$U���@f�	_��c ;��KSI0���v��g;�`0�^�G$~H�ezb�ʁ�����{_˅�D �g����3G|�XjDH^�L�S�;�Pt��2C���7&Z����P���K��������W��	�6�!7�i��,'��Բ����MV^���z�CH��;�ZS�a�uh��:'�ʷ.N��	��3~8I	<�qWj��ꃦ%652 ����+lۡD�_o��g�i�(��]�6$  ���HAĉ��ѭ���A�X��r�������!��`0
����1s���kI	��գ��e`�]Rσ�>��G��H$��匜w4` �˩f	�6.��2H���Jg��#�l���0X]�V�$¨P�L-n��A�Oq��{�;�$-G@}�����,����A�AZ��$�����5�B��s�o�Wb$�40M�Rg0��r`k���( h����!p`Hg�����S�$A��~���΍���V�X�0NMǰ���b�ǰ�d���RVD�Ƨ��	g��v_N���s�� ]�d�fV�G�gJ|�t1qr�Jm!�fVL9����j7�g9�l�$�#4�W/�ǈ�޼���q09�=.��#�镊,�|�����&�G깎�ֈ��W�.w��w7r{R��t��K,=_�_�VjwFR&�a4Xނ5�2�QO
>�.wAQ��\� ��Ї׻|�8M,|3@oVD�Z���j���4iKgb�����i%�[Vc�E�Z����z�˓��0���d�6�|��#Ŭ�c�tc[׬M�ǲ�j��Xr��r��_�~Co�a�����S��e��C��	5��؄�����_R�$��RX#��9��"=�2�q�݇�W
yi�N��0W��%M��Ut�!�2rz7��`ױ�o���V����ڄ��'0�X�csT~�3��R>r���ˑӡ<�5���2��<���9:�Q�Z�n��5uZ�������+�>�R�wi�b�_�5�C6�l{N��-7٪ݣ��:���i4wk���{�����u\RE��5�h��@!:rD������V�*�%�ۛf��n/,�S�=^��_�iO�D5���sh�\[���?��8#z'h�4��tE��!ڴL0�!UGk#@�.xc��iIˉ�VQu��2gK��]�l�)"�:��OjD���.��[�[�x���^�7Hn����4r�":UaI�}9�$gD+Ε�_D�B�F@���t���6��I�l;Sf� 5t��%��`q��p����b]�`�D֧�R9�v�*�t����)1i�D�.��o=+��/MX�WV9��|�Q�n<?�J�>A�c�.�N�B�sDY9��~�c��9��AX�kLYl܍�/�F�[��;��p�`����6ֱ����s+�~B9;�-6�����?��KH�U�Z��������؅xP%�����bN˿I�P/������	�[����L齅PS�����z�q�6(� ���D���������\���`�.�!�ȋ&��ۇ�5�7�)�a����{G��~:;��2���5|ḍV�}�o���P�Q�ĔB�Iꅯ��JQ���yl�38��O���5�.��l�5����<b���څ�[c#�>?��P�
s��ǍW���5$��p�?�cV�t�,�1:�����Q��XA=�e�麑��b��������O�K���G�_.}����8b5��藖(�+J��>���D�&�=^?�8�"���v��E��?/)/g$��"���lj�p�!*�#�w'��x9�����΂2�+oSJ� @b�q��TI�t=^�Z���#�y'�,������1�!3�����TTsZ�������cTݬ��d�A����r�7WA�C�S�v8���d&���Վ��ݷ����q�\� L�7j���^��-�ev��C�������z����1Cg6��1������WkZc��n|sa�@K���Y>��Aq�*��:s�Xe�����x�*m$y��X�g˞��<�r��]�!�8r[ڌ9 SK*�r{��?6�Mg����չ��\�P��Xq�ѽ�!�a�y\W����0����	�ޯo��]�'X��ao@�V�n �x����������X���&3حd���:�o�Dcn
��ki��0d=imŀ���G�	D9��)?"#A��ѹ�s
=�z6p�F�:�/��1�A��c:U�e_��	� �2��� �Y�H
@!c{C�ψ!B�c���M����G�f�`�P�}R�73�f��Dsh*i
����20J����ٕ���Ɇ�BK�I�xs��;�OPM��.���
� ���v��B��Co3M[���0>�㙤�u�ޞKM+��+��N� ��%&�V���W��n���s���섐�^"��	��&�Z�tf9���8��T<�>cm'���M���'b�Z@�'�ڛAR��vU�:���T���٘W�Uj/�x�r�Ŀ6r����Y�	W�
�?7ր�Ȼ5��������:ʘ�K�"��Ԇ�����8>����,���}�"^d�K���RC��ă<W�F�4�p&�i1�x�wS��2��A��)~����/�m]>�e��}�	��X�;�@� g���5��9�]X1$�A��y��� ����[�9%		$�Phi0e���G7�9J�����ԁ��1S�WiQ$���8�cjѲ%�a!wR,���E��1Iz��Q� ����
��%gl9��H�Q;�o��0ǽ+����N�vו��P���S�������lhzb?�X	��S0��)H�XN
8~�9�R��2�^��G1<s�c�/.DC���������c�9��BAb����`+בo��"�Y��Y��6is�t`��&ڢ ���n��+�j2ٶ(�3�¾t!�IK�WX|�@�dx�dvJ����v��f^.�ju�-`v�MEmN"T@�!޺��>O�x��ڵ���'ewŠAVF�75���d��g����Fb�%0>��f��(�~N�'w�u��o���ٝ:�h`1�ޢ �| �-�dAv�Aj��5�	�NZ.��7Bl4���e���tvbmQpf���ʈ 9N����	C��x~��&�9����n(���鶺����0+Rd[�D���k�����o�/�mJ�X�v�W�ZXFO����הw� z�eFZ���	;ĉ~M-��FSD5��q A�x�8�V
;�b	�"N@��)�糑���UH$�V.�:l�_�/��!�����n�Y�<�����
�p���p�w�JФy�V%t�ㄪp�]��2�A��A����#����m��|����y��;��"�B�d����匕ԑ'a�9}����0�jL.����(�+a�S�D�u6J�e��w�O��9�Y
Jےw��� �j��=�O
�]����O�6�F���3�}������i���Ҙ�{p���M*-U&'��N�q�orߩ.^��KS���$jI3���)XF�O����]]�e=�*��)�C`�-�C]�y�]@��JV$X,s69G�����ܢ��"��|��mz�[�`�H8�>���,�O~�$}���En_$�����"�.E�9��bJ<�:r'��Y����72DV��ۼ{�t'�m}*2�&l8,�ЌHUrW�e���	��T���byyj��i^�3���UpDO�?���L�R)���"���D��b����F��ǭ÷U!�����ΫX^�yQ�SKd֥�LN���jjf4�@n��ע��K#[�@1}�C��}G��eRճW#��x8>J�;ݽ&�fBt���V+�ϒ�\�M.��y����L�/�A��d�yJt�ݒ��G����؅jos���Q�|�ͺ�W�UcA����[���x}�z������6^����%h�<�� ���~X?|������jp��ܼ�ŪSbH`���3��xZr�o�*��{�>6�94�*��MF6~�>V�>[�[����~�g��;���@T���}-�v���?1((�y���g��M��e�y���~P놞|0b�����A�5V����_e��z���|�UG)�w��G(@r�id9�Ԇ+Ɣ�]f^7����1� L�8�M�b����b�|S��Uٯ�tY��5��1��L��\{~���N"@��m^���Z��c&�"���r4Ej^n8CI�/��� �+)X��2-dĖU�//�h�
6����L�%��A�޸���ycB')���&��+��r6���I:N?�PG��0�@S1Ho]�>�"ģ6�K{���B�Ƭb(��D��Z>�=@ G���V*:}����V�}a!�>~`�Y�sh�x*W�.�h����V��tN�8>�T�c��.軙"�m0�s�$�9^N���d�]J&Vfd�/|-Jdm�?Rfܭ��[�S����o�}N�f�`�Lm��ٶ"���@	�i�����s��!=XQA+�.�G��!x'
��������Ͱ{��fy��s������-���ce��R�6��~h�Z^����0l��k�)V.�C]��st,mew�Co�����%�M�t8iB<Ԫ}ì��Q������{�ȵ�
��MK�2�̑
�'u��epy�c:��v��ɔ��JK��4�)�G�kI���a�e��,_À��
�H!��%�@�T��vg���ag���$V+��0�q(�u�7cR��G8�/�9�eI���?a	��ߒ$!�,��iX�����D��o�/�������!~�i����J'/����c�Ǿ7�p�b��+>Uw���mǹqZ�$�C��o s�	���@cc�5�GT����u��S�5[�,!O��I���Hg ���~����%?2+�� �Py��_dW�L��6�zm�{�[�k��-�|�z=t����)r;;*ҾL
�4NH�H5�0:�+�|=���O}~Qh0��	հZ��<b�"���En2�aw�H�;E:�>��j�R	������A�'�&tMg��؃����y1�4��0�x\P�a�9�78�c�Ǭ��Q�E�i�9���c����HB�	,�+���e�m��F�V�,�#�����?�p�dA�\�}��i�ea����������,y6	)_]������؉[`b� ҁ�fq�9R�����oFU�� j�(`�T��Zqn�s��w>5�3߫��6z�c?*�q=�W�*��RY�դ�D]�à��b�)�p?��B�;ϦlF�4�A���s4a�^	=�̨S��s��e�=�%%>$X�1v�$~���k��;�A�����j�X�EA���#�'Ó��au�tw�*�T|:��P�@�����.��7�i�7�)�W�GI��Α�`E���ak/>�����^G�:��������
,%eӌ��[&2U1pO�|��F����B]�G]J?Қ*�4�$pa��'�b%�-dz^2��~U>��F��ʅO�H
Q}j"��y�c�@���.��LӦ�7����/�TV�0�M�}A%��?�t����9��X aW�s2Y@̣P��M����a��a�(���b)��bƫ���5�Ѫ��N���i�`9�)�V]�F��r����V��kCP�}��*�=����{�� �k��.��Ch�Qxjܽ�i�X3(k��w�wEcf����҉g���z���i��0e`��EfwV�㉃Br�D�@�?��d�XLJ�!��]�e,�������U�-�+|�ɑ͵Dr���	t�f�=#���w
��!�4�����*̌��}'�"�{��
���V@��!�K���s��9U9�h�W��a�'�Wv�E�ܑ-q�k��_�h����=�p�o(���~j?�OP�k!A����4%�5~gk�xE�0Nc�V�ؒW�28�2@>��S��ɈF�7�i�!����MpOo��!^�ǯE�Y!�)����-h�# &��񞙤0���R_J{��Y�0~8lݨ�=:��{t�,tɔ�W�TH
z�c��Yp�����.W ˅<9���p?O���o����P�\�\.�o*aU}J��.Z:>]
?E`�f��u:.2����c��ƫ>0��[_���c<���Y-� (��{L\T�����u��BJl�R�����$[�̽�tw�u��Ԧl�,�r @G~�Um��2���$��˵��̹!������0�jbk�/�b��*�!o�I	^�0G���]��3�F�#�TC܌�����E�^�d�
M^��6Xtu&��H��O
g�3�ߝV����)th6���ɜ^����{<�2����At����,�9	SiѦڤ"B�,�
�g	)1��`�l��r���+�\�G��lj��/��E6>�U�Sc�`�QKNx;r�J�ݹff���G�ЂU˻L�׭aL�G<��ތ�8I�Y(m�q6���*�
���жg�]��S��}� �	�^�$���_J�@�(] l>�a�땿�BL�^��.�J
>�7Y��4�w�6�7TH��F��5�9����=o�ѦZ:���vZ��Sȗ��W�x.4�M)G�N��2�6z�L�%G�E68C�JVa�=_��isA��3����^���L�9�QY���˱Z�׈�r^"`$����}B%_K��ã��-�i������8˸t��W�`Lަ9�G�-�Hx��%2������`$�+�x����H�.�X�����>��d��M�x>(� �.��k".�Y� I�85�F� �t���ؼw�� / K��K�R73�NWͅ�,���h��g��Yc
{FΩ,F���Ks������A�
��:E�?@Z<�P�Ip������B�<]�o�����Ѝ�2H *�=�{�9u����gK/y, x��E�$ �<�J��@�mz�px{-��)�|�D��I}*��-�(L(�ʦ^|{R�%k�ޢD�;�r<�fJ�ݥ�c^D��6�S�P�is�,�nJ�Q��}ޙ���*���s�3�����&*�l��1H��Y�$���gE��ʏ��_�|���b�����@����6E#^[U#��"9��j����P��j�B��p���bW��mP���G��M\��;Ӑgo�Y�jRYi� ���͉����|{g�6�y����&�G�v�ʄ�o��I^��2H��:��7Y�z$yvYD�F�4�+�������f�Z|��W���|u�咬�]�����h�d��hx�ٳש=k��4%�,����/S��)�%>�<��k��<9I��p��xAh	��q�c�+h-��*�-������t����h�K|�#^����(�	�Ai������3C��rZ��R�F��A����>$?p�H>���JG�׼c8���ӻ8����[��ޤ���u28�*<���G�~�(��#�)�-5�.б`E¸�Gh��i�z�R�"�C�e��T�TK�FC�����\#*�5��ۓpb�+���>� �ޗ�%�h �WR����
^䎿���A�78O��X�g:= ��	�5�(��-C)�x6
5����S��K,5����pAz�٬���J~�'��w��Z�����P]-��ڀ��u_�8B����To�1K���⢂���Y�Y�Ԭ��p��S�:��1��,C�z.^��^�[�qQ�J��i���G��>瘔���
���M�`�j�@��#X�w4�.���uN�/ ��'�p��9�_Q�r3����4�bxmg"р�R�
�y��֩ �8)�6�v&����G�N�4���:�Z�i4v���51l���:��>ع����&��-����!�mw~f�,�:�#J}E�S�x��Gg�m""�ˈΥtڗ���C]PzYC����ߍ0��HqO> ��5V�Wb�������J��3u$�y�>S������ *W\�ˆ�B��uvq��'sY8�]�X�����h���iF���>l�3��3���< s���[L��=re�+���Ė9p �O
v1bfΓ�`A5��2HOx�M�bzN���F+~�����*��A�-��)�sw2�8��2�����A��,�c���^Z�tĿ��������
�N'�H6Wz@����g�1> ���iM|���ſ��ha� GHK��z"1
��m��zΏ.#C��D���b�Ե�֬ø5JΗ���o�.ye�Z]6
����`����.�\rn���B�����,�.�gK�G�冴�t����g�+��O�s�J��)�P���M
^�Q��N�8M:�����^*�n��g�Զ���+��GAO(C;�z��;�^c����`��'"a3ᆋ���������������I�k@0���@k_|�����%�I���U&�n��_>Q���lU���{'����l�ל���0�A3U��cUĀf3|3Z��YK��B4G
HjxW�N�~���a���@�nB�WǢ�i:���d�6
lB���M��W"?��Md� A��`{�-eY��D!O���4^Z0s'TY��Y����|"�_G ���t�*	�mw眻�1����4i�7>	�L���Q�66G_� ݔU��_��wǄ��{,�ev���3J���z�F��c��(Y�DH���nV��r�q��L5�>����{s����;-
t�T�PaH��4U)?�x�߬�*K*eh���ҋ��Rg�͖Jj@N$׶����V�#���� ���n�:���u�ξ�3�r%������Y�jD�_B��������PW�鱣��\��y�?���;jß��^|��}�{'>��J�d!�Q��`i���$B"���G���B�Le��?�!$��"V�K����[��ʆh&>Y��_�@��ڢy��]��dO�݆��Y���.쏯4oRZ3���v����|'�E��p�h�iJhk(B�T�e���/̑�]p�'ۛX�<)��LC�i��$�G8����'S�P��uk'�ݧRHXL���0	n��B��2Lu�9V.�TM^3�%"��]�A��&��e��j�b�>)������Bk��T�Ҧ�ܤT'/��M�޹-�m�a\�kR�6��;|$G�*_�2wV�Xw��Q�_��'���LJ�Ŋ�}Ʀ���^�g��Zs�� �磅����.��E�$�c3���^d�-�Ѣ����H�h{��s`�����:!�\�I3�
��*�/0r 6`ƞ�$"�k���[8�P�U��;�7�1��F�R�u�8]I�_K�L�K�+�ҹ�}%'h)f�� t�,��� 2��x�]L*|M�i_�#>�� ��i�ֲ���x���hp�[�������`1�Wm�E�)>��0mL)�U��9���Wb���B�|�&��9n��"M���8a�ں��T�x@�W$2��+ڣo�w+J�5�m`դ=A��6v�8��$]3���}�G9&�)wk���4&(���c�#K�}w��H�.J]�&�u 	#+�J'=�=8mȞ5{�gɴ�<2�i���A2_�iù����H�����J��A$~�������ܤ�%�͎J���W�?�稀j�ȝf������*$�C)�Wz�ʹQ�Cwmy�S�W\�UV�}p���퓤٫���(p���T��c�s#g��Հݭ���a��{n�
��G����^}�jJ�mki�n� iu���+�e����됭���(Ug�����b���W�1�cn�x�o��O�rD��.�K(�l��'���,�m�0��LI���S5l��CH�����yA���߮y;l���ٗ�\]B������W������ˁ@.�I0)��m��lN����"�'��J�0���U��֝/�&@�F_K��o�LJ�h<�w+�0�D��^Y0��Xs'�)@"]M^�x�5����z�n�Hu2G"/ι�$�Q�8������m�O0!k�n!���UݿN[������ְ�*$U�5����2�m[��N��G��E�OJ���N6�䤕�k��^�$����-�`Ѧ�q<���Z,u1EF_���I�}!���І̸��H�X�BqZJ�������P G��7D����b�ɯ�4A�f^��F�A�&$.6kX#�7!�7�O0"T�1
LM:�e�m�'(`}����Ǘ�P��B�r����e�B.�k��M��������c5�\��Wֲ
�����:��S����r'�'�Gx+�0O����~�(LZcK�>z��:�`~�3ʾ!��D�*8XM�{ݺ�������h0_*mkJ�A�5��stK��`*)�H$�\� i_���G���+d�j[o����_�����<�=�����d��o*�+	SV�F���sU��A��A�;S	0�$_���M��]
���Aa�SPJ7A#@�FT��|�E���,��_@���mr�O9�qP��p$�6A\7R�	
yi�8�ic����N���$z^c�^U��P�Mi(�:�Q�)�#�yc�t��~	r�%�ܮ�����ߌ��t]�g��]�'�2�q��g)�e4��P?�3.<S����0X��"�D�,[+�#My��1��ĝ�:����TPݠq2�A�3�݇�f�Ϊ�DW1��x����ɘ��s5�څ�2��Bh��ަ�K����nXW�ұqvt.lZ�{'�r�M��DX���G������(��,깳Ї��T���h4VԉK�Υ��P�VeX}M��5;�<jwXfR$��#o����l�=�̄�=�x�^��8��������ٍES#َ����Q4,�=4=� ���+E0C8f��|ZA4*d/��E~:�x�;���G&g �	�-ɿ֜\Yp0$��`O�7���!2�\������ӿ3�a��i�U�����4�� SE�19yII�t�{�}-hږ�Q��e_Z��(����R5�;4g����� �m����DĎ����Y]-�5�y���	>��!{�ݿbb��Z�q'����Z�o�����4uی��e?J�Y�J]�XP�#F�8h�����Q����sn1�Y��R?�r�z3����R<�;aEMFϐ���1K�h��@;����}�ZZM���5G+�#W?�*i�!Q-շ�e!F�Z!���S���&���番��C�N���Xs�M=4)��K��_(Ϸ����ߛ �m�	�e�fB�X>��o��`�"H��f��6��(�H���K�j
���Oi=�F?ϡ���d����,��遟�X\9�0:�uԯ�x0������l�w�3���%�"��Q��`����l�v��w`�jp�;=o�cCX7gIy���C����*� ��:��:��Hv��Zb$Uxz��*��Q��|_<�+e@�e�e.C-�ȗ��3=	y̪�,?d/����|X_�MC�Om�����Қތ�Y�v�-�}�h�긓�$��rYs��6K"�Ap �[���"���9ה�D ���j؉�e��xaP�t�K�x��.Þ����b�"������yiB7gd�mxA.�#
�D-TI���8#�I�$��s��8_1��O��
M�����<YH����?qr����>��/��A��j���&��l�Z<�M����0�G�.���Wg'���d�w����΄�$��j��r�`�Y�0ˈa"��i��_��O���!+Q��+L�~G����p (�P2
��ƳpG! (�p~j��Kx�:��ٽ�*P	�3м�8{�>���)�����p�F���=��0�"�8A볶Ҡ�Pmv7z�ū��ƍZ� ]�j��k�7�D�7.��D6?���?�ύ�r��v-��3���^��9mI@��{������cƜ=���Vږ��̔�#٭0Ǩu��ft�^���du6��E�.m�[�*�pnCx���."\k%Z28�綠g�a��7Q�6#�|�b�0,m:iĔ�t� �`C��n��Oh�G�?�}�h\p2�i�`��c��xAP��n0{n�.%;t���8\E:�A����~��c�-�0͊�ī��6M A��p��n��6��>eD�wl_F?������ϻ*)cF	d�_�8H.��J��������EʯB��0��%��AŁI�R>�I�Y��b`����Ď�I�޺ʧP�4�_=9*\��-��P���?�˩!�O�q���/�-
���u[����I�z��?�_Ǉ���0oY7C��.sl�8��{����Ƽ�.m��:f2֊��/���pv�q�3�r)8��a�M�Y�8�O�:��+șw��f�}��JE � �_?�����D���
�/�Δ ��������+����ݝ+=�B^fi&�f�Y����_-m	�c����@,IcCa
	u8��5|�a��6��{��n���Vpa3s�~��tU^^��U�-����Y��	��<��q:�C�"x)��#дLd#4k�Zg�	��.�2S����G3�U�iO��(5�	�Vf��ʠ��k��ָ`P�{�Pu}���\n8:����v|����S�!!�&:G�?�C?$y9�%�>��w�J򁗑p9x�r:�데��:���3a�]�1�V}Y��)4V�Α�^�*p� �!��k@���:��u�6,�`E��^�OSG7[t)P�y�F��&F��Ώ�:�s����<�b�lM�7T�Ժ�`����m֒û�ty;��'�q�y�l��E��0T�q~����X[���UH��(	�5ۯ#�BBbpn�(N�K��/u��%�y�x͐�B�� ]��h�y�$=ԇ���U$�l�*��jf��������M�X����c`�?Uۼ��Î�ʓ'B 8���Nƛ�:>�}o�☫��:�S�_��Z�;{.��xO2=�^�K���9�Ù����Or�@6��J�FۦnGjKK��t9c�m�foWt˝oN��m!��>��!���m�r���ML���@?����/	�P��tb^p
'��~��a
�qId¢*�A)��7�'�������@�W�Dۂ��D�������}�}����`n��1G}(�@�9o�����W�p4tm���y*�¢�v�wee�(�t;q�d���#)�Y���4���m��q(E��=9�
3��.'-�#/����)R�8h�f>X	N��3kVJsm�M�y�6qW���<���\�4���yxsσQ��Uɷp�4�&���׈^V�Y�(|r�m�F���8��Y�`�d5��D;a�L}�	�|P� Z :vC2�ߟ���f� Xo����Fy��Cq��R ْ�ر�L���6��-���O ��,Fy�{Z��3�wrc!�)C��;Y�$��14�pGǄ!l!����!�#����Gv�8&��T�h�mC�t�MfzNή˨�i���-<����e���8��Hś%�H�>/1��P��;��5��A�t"�J���2(_�lD��>%F�g})g#|S��,�t�s�`��V�U9��)#�Ϛ����K�Ϭ܆\�B�5n�0[��zذ�,C?�������G�a=�,���DB�r	]�}�/�F���2�o���Me��jh�ȼ��<�Vd�R�rX���'(������)�v2��W��w���_������9Z'ɇ�����Et��*�G�5o�_� �]N��Z�����ҳ�ƪ����O����rZ�iCR�͇>n빧z���ʣ�;�#��p�y�7���hW1[Oi��w�Nu�2l/ sQ\�q{��p.�;�d��$�/(t��u{�E���1��MRu#��gOô~j��!�o�_Ξ�/!��	����>�f�١�T=�϶�����: V��CW�vk���\�x^��oj���ݪ��D����|��:t�%<$�Y��@�8(�� N�{։%Σ*�c�=˨�磔 �5^b�~�0��+�a�m�7 ���� |�7�]k�m���+��b 9�?�b���[Ņ��5UyL���k�_Y����A�_x�'��;�s'��a�"�Ҡ�U:fWB(�6r�c"}9p������8\�@��~�-A(Ϋ�WH���	8
��ڒIgQ҃'�x
�'�5�T�EѤ*�$ާ�֖�-v���G�e�9� ����gG��n�$(dW.bo� w�FԎ}�|�+|`3}�p$�6��d��S�ԧQ���B���Jq�������B�)̹�z��ݑ���G.#��p�N�G&'?�[3A��XP�H���Y�/�b��3=r蝏0�h��WY�t�m�Xȡe]��^�!�4�vx��"�i�S�R�/;�[y�E�a�-[c���|�U���=&�g��*�Ai�FA=�zx��.`�n _�Ŵk��N�0��ɒ�4Ιĥ�ee�v�8�JW���;ϋr�`g�>�4���#@�R���:T����^��[��e8�<�
ʨ�vgeČ���l�LqJ	��s�¥�D��_�K��3��J��%���P�����L�uN�m���.۱��]�M5苂���w���1��w��1Dxf��P��Y�~�����I���Sbǡ�xt`:���o��&+�i����J���>g��F��Y����VѰ�{���6�'�<��`����>9�h��n��>WI	��iu��I�#ǅ#�d���-�VJ��E�H���W�kU�1�j�̪6��X]�v}��Nζ��s�9	�b0�?��:�=�R�-uvm��O��<3/n<�g*�,�/��c=.�Cz�y��ۄ_K?����3!�m�Ui�b�=V@rs^�A2|~褷�*^�I�M,C� ��a�.�|�cp�Ḁ�9���G�H�ʄ���������0H��uV�
s���C�QWjߒ�I��mE��ʓ�d��l�8�q/�?0��-�e��y<��>�l�z�=ܛ~adg�S�B[W{��^-z�$)��$��T���:vaś�c�91��J��[_�<i�O�
{s>��2њ�XWՔ���D�:�M�b#aĀ��r��.½*���J�F�c#��
 ��zV�0����3�x�:I-u1�|��|�P�\�$F�j^���K��W��q3q�*t��'���dS���gw3{(��	��H�AѤ�`N������ZQ�@�����,�4�D���#�������� э�������ttdeql�Tpq+�P'D���K�+����c G�MA��6�#p��l��<�B�%%X��D�ƍOOo���>I����D��u�Y�}�~ _�X�W��Uwj"�Z5%&�0)��̘�~�(�<x��mKbh���ib�B�4��,:�T��cT��joߢ�$�A�x0=����'��Rm��&t���:��u�ß�S�q��%u�vEh�ee�	�T�k�ʦ�#;�,�<��ZJAH���9�ې���Š_$CoD�6\>Sjh=�>%̖^k�6�7����F��L)�[���q���L(2Ocy۸��J|̽lz!��X��#Į��B�#�.�J���`�@ot򞻳��+t��.Йi ��3q�7#d����������:��Q�`�x&�3�H["��br�RQ��ۃ��zG�^S��v��	�)�V��W$C��r��i���|����ec)��ByX��zp����帜13���+����"SL;ۖ���S��Iq���%g
��C�̖���\��?)���J�1�H�o鸦�A��&�Vr�D�B�����޶7��l�o����p��#^^ɺJ(Q���\UL��{�4{pz�����'GD��){e�Š
5�	�0�K���&�����\ 1�-ǧUâ�p� ���΁�m<eh�»�~��ԏ����&��9��# �)�*�����`r��B���dc���}<P6e=����D�.J�������ؙ��e�N�����3�:W�)2T�r �[iG��"�@)�	�To����+���:���,r$�e:0ry�\��F�~sc��A�evf� h�;ui��n�4|ǳ��Lr�������0���P�6�/�OO��.�'l��I�%Qw�̆G4����[�+�����+.dn�"��_�'��$�Q�pR��A�a�P� ��JxP�V���������!+n��fs�7ZQ؄���჋�'΄oU:o�'{x/I ���Y�MNXQ��S�dY�� g'R�u��i/�S���Z"U���J⃇3�J0�m��ʣ����]bvf��σ�&\�ZF�G�!���|˜�B\Ww�J�Z��F3�a��=�c����	H�`���C�Τ���b���C��ĳ��M��E4R����@�a*1:e��;c]��qO�� I�@)���[��$4cԥ:V=�L���M:j�u�/O:K����5���J9n��m!m�O!�I�{�-F�iQ�"����Y��^����`��|�sz��X_O�5~<\~���F��c��Qm\�ح�K\pIz�$^�u�R�� ��x���j�A�j��\���o�ģ�3�
�Q�@B���
�V��ݠ�v�iN��S�N�F(�{���u��B�|�Y���3��o�������亼�M�ߜb�٢O��(�2ԋ�43���_4��{��m��~% E��a�Ϊ+���T��3�g`���֩kusI�1y�������i�
�
��m�5
���/�Q��R��
EJ#�)A���
��mdS���E��VKg�['�z������F낕E	�N����t�8�����Q��y�k$ �U#����������4�p�t<�����ww��m��Y�����?c����/�I|����\�����#�V[  �A ��3���1�5�ݯ�.u��R�ㄤ�
yo����?i�0#�2�D������U����k���^�׳�>�����غ�!��>�H�4m�q?JS�������f	��`��$���[r�����gzټ�5ʛ3cJzIn��sf�o7�<���]����r��\G�:�4V�;d<���%|��Ł:�5���������{�������b$ډp'g��
�oL+m�Bg��n�R�Z�$���u!~t1��o>\Y�3����0�Ӡj��=B�G��}x�C{>#\lB-]F<�X4�1@R�s��U_p��kg���aƯ�0�鱕��Ey�C�~�\o��(3�C/�:�aN_���=�L�Ò���k��ȝ����7]�n.���3���]<Z��qȸ�m1[k\������P�>=��k�����?f���z��"hn�7^��I$��@C��I�ZR���������C���@�^�.�>4_i̀y����`��v���z�/�UXp�<�el���V�,p)�@C�p"�ȃ�"ke�2�r8ȩ.��?�x�x|%�Q.�@�}�";����B�4Y��m�୯	�܋��H]����­�J�$����Q��S)l���� K'%���OX�P�T�~7+!*�,і��rCK�e���M}	��K�<k��
�>MN6F�S�@�Z�[��C<{���x�����"|��c;��7 �iV�����������o^�?��*%����b��h.�?;���!�p�s��^zI�4 /�:!?Ȱi6�o(r6\絋�ߑ��%�r�E�����c�yh[��Ͻ�͇+$,	�����]#��jm�٬��ظ�AD�L��Q �P�1�{i��/>������P�3��K�z�S"=-V��>cL��[��:�0͓N�vL;eg�;&�J"�j�Ѫ� $����N�n�&�z�T �U˖	�q����{1	c@.Dy�o��ĥ3ے|x���NY���<FƠ��ܖ��}2ȝbx�	�8R
 �ͽc�t������*N��>A4�2S�G�M���W��5����!��`�������+K?���?c�&�}��Oy����x��.���� V��Młs|��s����:|��x�Y`'�U>%�F�?�t�y>ćxJ }\�$���P��SP|�.�=�pMb�	����?��'n�sJ���D��������Rt������h�B@Z�c%�
Lb��I�5Y�g��JQ�)d%4��&4�jP�P�
n��erlC�������|w&�H�]o��R�H@=l�Y�RV�Zѱ�l�`L�v��<�����x1�� �++�|������7:Uq����hU�R å�)�6&��dh@i�L8�dz�ԽiU(!}�3���":����r�n�����z�v�,m�X�݇�pOܞ�����-e=�(�𶶃'M��-�J��U�ڍ؊���{���l8*�����ūm����<��|*�� W!W0��z&/ҊuZ�����~,&P�b��@]�A
��8�C O�]0ɸ'��������A+A���],7��KZ�F@Z&N��:�Zl��P#�:8[~K���=6�2��u�9є�T	*AS�T�ƃ�!����N/Y���3^h�'��.���|����cX˪�8�d_��!񐵐��`��|O T!L=�I�����L��`{��r��}�q�;&Srr�MoA�^ͅ,��?����?��������Lp-�Sg��5�f`�c�O���`���F?���HȾ�u���=f-�m�X�#���Kj�3a�Hq2U?w0d�9,�j���,ӒQ�*�M�4��=���Rxr9t�g��-�38�0�U����YU��@Y��f{�SR�B�X��t����>�8kP9!�_�1�,�q��lPS�L԰^�~���1����{)��o�V+)�(�3Ӊ��]�[�B귈㋸F�@�T�WR���恭ݥ�bڎ��w�Hp�\����S��־y	*
�)�}kug��e�H56��,a�c4�U�#�AX���f�+������5t!��I1�ĺB��૸^(�G�`m�;;Gݮo^@�a
���
O@%k�5��(�T�6ȗV�a!�9��x��k�P�% �Y=gyG>M�,��qc�g��K�g)3����u�UF|q%�m��蚧���Yv����l)D v�wCa��%���T5-��l��c��s_���]��;�-U<qg{,{�������l�V�7u��)ځ��vƧ]�".�fd���������ǖqu���>ЪrU�iA26��F(V���'h��g�o�Cn����oB7żN垅|��*d$�&���� Uǝesb�d)�6{�����0 U [���%��l.�:�{S�?Ě���Q���n��t����Y���)��"�Y�	~�_#\�V��s�7�Z��v�`��l��J���p -�!Ŷ���P������t�rٰD�:���r�r��Ѿ?����}q���A1Ti<	[�h���e���|�2��E3�j��e�l̷v��v09$�̑���=�q�y'9Bf7�']�l�*�Bfd���er�v+����d[t�X�`����Ѣݢ���"&�0HRecBۇx��ʟ�𪭠�F�>�ݨ���&?i�@���rG9J�H�)�g9Q֚���bcM�e��&��t
��
`E���U�3"#���<��c?���Y���|W� G����Ƕ�[z�|��M�aCc.�������#���Ln����=�A>�@��Y:���$����2��2�	�N��2V�X������ǖ���zj�&�I���)�(��1 '/��1hr�� �%��E�v`P��[A�7tW�|a�U��F:��] �b����ד̳[{�������a�Iݨz�#赥��TZ��۱��v?z��$!���R�I�ߔ&#�!S��Qe�y$0�� 	C��(���s�
�i�Aa�P�*f�?�z	�~N�͈�ZT��]{b����7sgם]�P�����k�%8z�����J+��y%��.����BLm!���à���*�3[A+K���}l�y0�$�/Mpj쬦�Ժ[�*�f��X���+l�@M��Vm��� ��mrN#3*��x���"Q�K1�2" P���g<��V�L&=Eϖ-�g�c9DZ%es�X3���eV�!��T��1QH$��ZB v��D�+I���b���6�'e�b��rd���������R�)���w�$��S�/]n��aGLs�Ӟ@qk���<��|q�p��xR���QFcnq�]��+�]I�5Cz���32ɉ��r@�h�[�U��+��G�;�2�&�����e��H�6�({w2�9W�V����S@0�ľzcH����k��h�拤�&i� ���kc-�*y�կ�j�i��Zk"ޱp)h}Ueՙ���KII��c��%�
S�+"z�}�M#�b�`�ڧ����2�X�3����NO+�S뱦�&�n��aD�HA��d�A$8��4S��%!R����Ht;����a)F�<F�ؚFf1����h��i�ZS�8��j?v_
�[�p �Aie�I�A�����&rޓ/���}n�gD�~���5:aX����D�z�c;hk�(�֏����۬���xFY;�z ax^�_�;!�e����Z�vzȑ@Lh�`V��㪃 ��������m�9�vE@�.#���'\�}��x�#Wb�#����=v�h<Gi`>i8#v��������
@�|�n�pJ)	��n>�F���e����N/:B���B�#�'▀-�T�b���
�����X���p�Pc�'�X_w5<�ݾR`����?��@ం�x�sdŌ�}�ِ##O	*'S���wJ��ۭen���܃4�jm�4&9��e�o��maĨ6��Rp���f��)K��J>~^}п�Ξ��-{<4
��ڊӺ�s�?q	v��xs­��U�D����򂑓W�fX�^�8k�ZHɴ��&/�`$��s^G��%� �h��m��I�O��ͯ��Y`O��h�8	γ�$��v���Y���#�����0�|��XT��/
���Ĕ-&d1�Zf��ު��"�iJu�qI>�v��h)0:M��t��G�+�x�~|u��c6)O����l��c(M���pCQ��' �hin��͊���F,X2>�2wz�=�kh[�BlR=U���?.>Y�Sڸܳ�`SLC(��6��Ol�N�O�+!��m�c����2+T��xü�G㪦�_{V�������!��)3���vv:�U!-t�!�z�K��6��Y�4ܦ���r�j$�o����j���zK~u��/93�RO�(��L�H\�=���P5)�IM�z:o1�FSUn��"c�u���:�xU3SRR���R�dU�Wv^���k�$`#�U��8������$C���`��"�{��Q�ZS��?�r�C!I��g"/��߹�؍�[b-�Y�j`q-��*k��
��M!�ߊv:�Z�3���u����E
������!�)�قI�Lż�J �M+!�G����6>/������,�o�r�^-=`h��Զ. �M�k��3˶J��U8 ��)�:�.3If���z�2d��](c�����R�>����Q�f|��٢�{]�ѕ�Nv25AJ���'� y���;��/����'6�
o�񣧳�m���q���|������ǹ�|�G��"�氊,������k��@$r����f���ч���Aq�B��-�]R����ĩ�ܾ#�qr��<`	a�'|q5�`Dś(g�%�6���YC�j�EwX3���HK=7�*,r�Ku����(dg���YW�|3a�Wዼ�B�61:nt�-���*�b"}����M����D��6���>�@r���g�!�7����p�$̺s�qA.����5n���D��l�%�N�b��̠^��O���
�"�C��/�R2xu��+�$���|,ć0�Yz�SLohH&��̭v��]	'	���R0�3r��/�6���d#!��w��0U\�g�[�Ǭ�B#9�"P.ؾ��]G�X�ĭ<1t*���'�|��`>E	���''Q�VOՏp2��������	��q*�`��r�� B���2_iu�uY��t���e4��K��ITjkԛ�f���|���L-��=�S��1��D�rH�u��\�<<G����J��n�ޘ��?^��@OB��L�[&�����㴹�Y {��"(�曮�Gp	���J���pp�`*�5�Єw:��g���mh/���(GU����x�A ��Hщ'L�I�s��dz�пK��X�Dq�I�}1	��@r�#�Y�A�������=9�
;s��������_v�\x�4B?x*�)���Q��B�����s�%��h����J��߅eZ�"k�,�9��֤����|K��>9�e�v�wL�j���.@4�Y����$��̩d�Z��'�O�x|
d3%PP��c3]���(�M��{�?IjN��pgz#D��&��_/�`��$���=�(i���U�m��2I���������0����`q�jKv�\6>�;tx0Bv �,�.�����_�s�*�����Aٚ"ml|^�^i�h0��͠��8��Bn����Ѩ�=�D
�,��e͝�h)b0�NI*R��
J�s��3H���ɕu���Ӓ���vh2J��9�P�J�	͢R��A}T�zJӪI]�w����m��c�p�G�Q����J]��&i��|@4<$._�p 3����۳}y��iV`PI!w�rP��K��I���)4�INS�.��e���E���DCD���[��'�i���`�cݎ
�o,�ժ�U9���ؾ��T]"[�����D=^��B^rj�6/��B�$���#�R@�'��]Lh]E�R�ŧ /��������Yb!/�o�o��*~���g�N�@�k��[v�"�����vAX�T@�~>���3���8�U����tοоw�:V~Bq��`�6�ϭX��J�Z-����=�O����$��4o��ͨR��凋��}�c�d���Rm�)�*���m(��I�	p����I_�%a��Nz`�qW���"Kw�G��v����1)lN�噖+��]In!>i�|'��z��{A�<��i������U���Pӯ��T�R��!��񑏋r-���dc�R'2��/���[k2D�ޖ�#�^�d�- swX�Y��?�4���݈�7Û�j����Q��F�!��,��@1�W��n#���*��B���n�C�G7a=�X���(o��������ǰJ���Y�չB��7SFQP��\��RgM8��/*��9P:����1Tp���AG
l�#��*c_Æq=�Ci�F�h���yK��-���Y�;nZt
N9�]�47��͚�<1^��y��I9ԫ���7��"k�wq ؋���4%Ux���I�j�������1�i���T�f~�%�E���m�q�����p0%(r���#&����Y�-�7��-q���#6�K��-���o����B���X�G�V6�o�]m>b�]�'�(�Zk��~l�[W�Φ7W��`��V��4�՚Aݹ� �Ro\���k/���;��H����b�6!�͊@�>�@p�`K����Spr�f4(ڼd_���6�{�$���ӴB��I��<�Q�S"`�n��ӿ�>�egA�4L@Q��`�\��vz�m�%������1�h�NM���3 ����I:�/��4�Իުֳ��3�Ϻ3��.��:�a�g��L3�e�<�s�?J��p�����<B����=�5>�M��2�\1ڧF�4�X��>��L�_����w���7� �m��of����H��K"���̞�L��t�4���=X�[+������8(F8��Zl.ߤ�nΕ�&C�H"[(n���������Z'����s
hit"m���<ݙo	�a[w�-iS��D�܅ܙ4�c_������>T'��Ǧ�S�<>C�oBy�š<c����hz`T�}�F(���b�3n:�ab�c��g0������ [oVw˳֍\'J+D�����i9˞d���烠�]~��	��M/��7�4���ȒD��ӍGV�tD��0%:鿻���S�����Z�5$���g�f��#r"�V�i>e�����`�j���
�=��s�	����0��,�'�IP$�glʃt���W�Wa�p���_��U7�]�^��3<�4{��=�3׾�Z�(;*2}��T��H/Lo;�v&j(�,��ץnM����Xp�9��[�����`N*/�5������N���V��j]PqD��2��J�̝�G;wk��S�?�P�"T8Q�(�~�с��5��b1�/�Ds���I�!Cv�fk��L�͏�H��� ����[# ��x��P��E�D�O���Ռ y�/���ms��,KsGT�_��Eo-�-��?5��/�]76'��R��á�
R|$�f�WN�� ^�D�p��BF�/U����R�nP�wP�xo?%��G�9�N�S'�|'�3��C�r�؎i&��*��7o9��y����m[��$�R�m��"������/��s���A��<B�\��L�ˌ'��	�'�@X����Hf�nh�a�rg�+��Osk�R= �s,T	w�\@0��8$|���E�_.�]�V*(�R�ۆ���	��K�~��t ӈ��Hh�NVɰ��(5u���i8�eH�:�p��w5e'�~�zJ�E\ĵm��'.?��!2������dѿ�a�>(r��F2�s�"��#�q���	�~�����+t�;���y?w3���9��g����˹C�T� kwglk�[R8/bQ�M?����5�rq����,�S�=�3��5$Ѷ��
�<TrP���l�tv����f]*���lQ�����0�`8��|k�3LHl~��lC�b�@�$*|���� p0,B�nԯ=�U����
�J��o �I܅'�jƽ"�=x����M�'|�YSX(�k����
��v0G�*$��V�����%�h~��ib�v��O�RC0��~�=*��?�����֪BQE���Q��]�z{	��,kD�e��GD����C"�ƀDФ�dCS?N뼞;��X|�{ߞ1dt�_�^�,n`
��ow���h�1�Ǥ�,m����R���Gw�D�rOo`�E�xu{������SO�Eͷ�u!2Х�r���{"��'�7ۂGeM�!���JY)�Z*�*]�L����$�;���#��wq4� E�J	�My�#��w$`#7*]�E^���떅nO|��e�B)�`�3�-����D{�y@9b��¦Ԣ�Z(���?�9B%���s�� ��ez����?�[ �\�=��K�t'G��bc�8�6�!Z��sS�* 8o�\�Ph
�����8���V+�{��K`
8�>���̚��9\wXQ��	b�`�d����c�Zx�\�7hX�Ha}�KZJ���fJ[��Bbg<������?_��R�I���F���؇�j�i�$���$
��Y2�h!|�'G�1�¼p6>hW�a�D���1�{"���%I���$����FoI �fρ�&�j\���W���0Ǜk��?�	E.�p�0A��S�v���t�c�G�P��W�9�-*�Y^�SO�L�Q�9��=�S"Y�}[B�1${.P�gݵ�d~�7�������(C�i -A�w����x]8p���v2�4�/Ŷ���c|�,,�{kQ�y���'�c��H����J&��8KDbQ���`5�bl�x�y���\��e�N���k�'�Є����q��PZ3a�{�R+��Y�	L֏_����Rn�1<\�ɶj�])j��h�Ǣ@��M�;�+Fp�\�+��!�mL�񒫯�K�;�e����;�T����x,i��������c? ����'�g�፬ ���3NB��I�k��6��{w�!ޯD'��3ƻ-��VmڷW<�W�(S�V����e�,���7�I�,�S;�L"/?
�O�cu�ȹC\�|>��� �t�t���N�ME�M�<7�; m�]�U���3��E�%�I'�p�n�=�3��)����I wx�R`�E��K���z���$m3Fb"�C9�i9�RՎ�����]S���=
�63$��Ne��C���8e�a,���XW��Ld���p�t#�Ϯ��m4	#�U��Tz8�r:O����>�$a3�[��H�f-]Rz�X�*��A����'+fDd5��O̎zq�E���n�M���&��
���NVɎ�d����͖�]�y��I9������0����T��Zb�V�̋����v#��غ�NL�q>��ӥ��4L.!�z�X=�:��8�f���0v�K@��ٻ[|���:�7K4'�@���w4
` P��Vs`�2���f˥/�@�"zM��TJ���o�F����Ąz�+u�:љ+�kJ8�`�w;�
~P�h����<�u�E������������e��<Lp���	�;9�>�K���]�~�w���JA�9m�xdd��K��u䪆n@o��T�/�#��m��!{�����"�w0b�*��,�7��=�R	�� )�N���Ԕ0�|�`���^��������X�Ɨm2hc"��ZX��0����ô�"�5�H�v�mu���2tm�s�iG;x��]N�>�ݖ�WI��n�;8Q���F�nH$*�����u7��i��	�~P-��v)�S�1���"�C���ӓA�U��* x�ME8��'�Y��Ÿ�[�b��uwgmH'A���ŵz`����C�vj���GWN��)8�ߍ� m�g&��� :MgEbW���n��z�́]�HT�i���;��m,�<��P��JN�d�g�f�k��l�Z�p%.����`�	�Df��h�����諦�D�#AӜ-%���p6��k��唦c|w�(�A%Fѡwue����%1N%w�X4���!�٢���KX��fLw��Ҷ��~|u��a�%�Te����M�}���rzBP;"0x���X���L��5�0��H7vⰍ$'&��A�'�����:!l�ʔGH���$vA5���kG�t},t^�co$������[?I�đ����%o�*�rZ߿	���w���@��f̡��/��s�3���I��p,3ڻ�CR�f���',KŬ	�|6�B�)E1�iˆ%����\�Gz�s
Z�|�a�r��<ڋ).���R�7W��	{��_pNDm�v�.G\S�;���Sѝ�%}7��Z�A��q�QC��a褁tD��~6����8���v�����wѝ���/���|nd+{z���n6wnO�'��Uh��KK�O��N
�3���n�A\�Zi��.U����X�����uF�cR,���x��C��G��D�x���t
�q�HO��ʷj�����q<����\f!K�IN��Gn��,���@��|cLw0
6k��'$?�k� ���8(�#H�S����bX����fo�B(�7�Ui�E��<��t�|�L]����t�A}�6ހ��& 3��]���|ۜ��9�b(=�اWCM�#H�q��v�U=�9Ή�̝ݭC�����_[���=*ֹ�u�҇����!���
�1 �b��o֢�2U!���%1�#A�����9���!��2��a��֡��w�����Y���)]�wI�E%L��J=�����q����%�5�|�����;����eS�]�7ץ��q�l�#�ZPn��GG�c�7,z(�����t��-�A�Y�:�Δx�T����ށz*��֦���lP{�A�i7	KHw����>�,h������Wn��u�����lxLG��Y܌�[8ul��Dt��.��@W�]����K�K�ˍ�cOb��hc��נ�>:�K��������7�6 2�������>v�=��K_Fב�*lB�*2�zu|z���48J�;,nF�e	�_�ި�Vo�1x�gf�s^����{�T���_�ʚ8+��o*�߯{[���/`�����A^ܰN�� �|����^'f�$�ITlE���,�{rk��d	eȕp���?8Iup�[ו'q���g9I^깜�
g�9��y�'>�}�?�%d۲�Ko ��їR#�_6�y������sD���)���E緻}Ƣ�<�IP���@��;d*�Q,(�-\�[p�J�0m�����g������u�n����&���ui��#-I�%�LA�o��Ƙ��c):6�smFCM�=���2�t�j��U��Ĵ��<\o�,�8o��6��d �,�3�񁲁��ۄQy�r��y%�����Y	��
���7�{��(�׫/�~�|��-����S��Z�k�����=SC��FQ��}ؑ�/W���K����E����v!�Am�f@6m��g�uN�U���^3\Z����g!82sՎ�4F|	�Z�^dQp�I�A�	0)�Lj��I�X��H^�CD<�}uc�h&6g���(N�+��
km�*�4�E30����'f���\	� ��$��q���k��4$_C��g��8�مex_��ș��Q�ٙYq���N�Q�C��-�;�~P��[�g�[�>�~z]϶{���h2K1�}<g�&�����q��r4�Pp�eK�p_�R@N�?@i�EԡUONUu{� ;g��=�2�y�BĐ�A��^C�+�E�`�-�������T&�q�C�~
۾E2� S��j�s���'E���# ��W��\&�]k{��e@.�n�Z��/�����,֦��	qq�v��c�%��/z7��^3��T `s=e�_[� �����VI_??'$��	�&+�F{cƲ�r�䅤�n�z�)lF��i�g�����N�%��^es������ό���iIA�Y���x�]w��T��g	M��Ա\G7`	 	��_���fܻc��O�(t1������_�a[�.�FN4R�[U9m�ِ���'���b`]�{/AU�N����f����Hܣ�a$���v�čl���z�n���N�^�@��n�t�wY*�!�49+��O?X*��N�:?�nʵK��q�+Zd��؜n�ގ����Gqa>T{�1��R=�AxU>u�	o�6'��9#D�80L%rqǐ�@�/E���R�$_��:�#�pk@e.�8��@��#��,�Cd"U��%c���9��	W[��W�~Zp.5�S��Ʌ�>\��ɛ��\����9��(�5��l��U	�� _$�V%5�'p��q���*1��iݱ7�;�F�D���h�3�#��*@/É(d��*�?�X�&�M�m���B���E���\���Ψ�̜��)9�m]��;�a^�H�^��|�Oe��Qrz�7��teg�*i}jc��t�x#�թ�w�MR�mġ_������%m�к��i7���!迯�N�56SG��w+��p}�[CW}�"�.���^z|>Z��uA!ڔ�S��t��x9���O(
�Q-��PU��Aa�����k��ߍm2�MQJ��Y%���M�'L�����z��bb�E�D6������+?���x��:Um��/�VSq���׍8��;-��\�U�� �����o������>��F8���`���G!(�)��I��}��e�y���|)�d? kE�*��ُ�����e*<�$L����s5E��/n���=�Y�!}A��mx�4��:N�u��@*��8ɏ+�p�@�����$�l�!qx5@PaF?`�U�'?��mP���01�MZ�[Z	.sd	��#QFfԆ0;�4h�D�y��*�������<5;���:(�[���96�e��xW���Y`a�慷⦢�l^U?>"`\�������z-�����.��^��3��h��vm��-r޿a���T��v�: Į�s �/
�=�}
w=��TXqJ�2��P�^�eK\��-%6��#τ9�|U�J_n�㰋%A��_�Q^�殿z֨�F��8~��c���"n5�G�ɷZ\wO�nȇ�sR^{��l|Yo�
q��h^��p�ʹŇZ��{ˠE�������:c��ht�	y��,yY's��od>����%�Q�.u
���ѝ�fլ��X���s��K�jS���%8��4 ��xQdr�zb�kÔ���H۰df�-�*�E8>//�J�z�&u؊�p$���nM���� D$8+[�սuxCGJ�b�.�^A����9��nw~G0��Y̊�E$r����r�Ӭ�H}�y�����کa_�D1����0������4=&�}'�^��:۠�`l��1�w��G��vu��҆������2?aK�gycF�17���Q��9=� �,LDN��l5�����7xM�N|ѻ����HHw&|���HD��5���t���+l���&_���"k|r]Z*TK��*+�p��4��(O:5�lz4���L�U`G�܊$�j�7�҃�`�^�v�L��׎�� Z��!����̦��?��;�h[�o�F�I-�Q�p�M��G���%F�A�{6�� ?��Fw �����l�t4�aM8Ρ�^`tۢ�������c{B��[g����☊q�{3",?vin4����:i�!�YE|Rn�G�'� I�}��r��˕F�.EZ�-��G�aJ��ok�nv!?���Pla�H�{9ٍ8��p�4��xj�5��H��s�B �ܺ魬�t��ۤNxwV"�k<����<�Gy�a�vU�]&V�����k=�IO��.7�� ;�֣o��zA)�n}U����01�x��u��wqW���/>Y�=���.��<���5�8��wR�T)����I]#E����h��rD6�z�M�Ȅ�CS��h�C�U�/�T���|u��!����l���IPh�Fh�"�� ��*n�;�6�&6K������'9;�4H����K�
w�O�!��$�!X�y<���z�.��Y�9�A��d���-� n�`ݦ q�����=��0�����V;�kD�>Ԭ[��OɅ=cLD��Ɇ�>`�H_����*�ux��I�x�@^N�L�53O>�lގ���桺�eA��Y�o=K��|^��Gٵ-Q���2�7{�gb}�?�c�{�7nm����䨼:�@mzl1�Y�!Ԋ���z3���`	��=�"sg�R$��\�m(�Y0Cګ�����ɞi��<V����e8̜Y�:��E�Ȏ����H"��^�J?0����q'�Y�l�_\TOB���y3�
As��.?��\V��")���e��|�����4�]�:&s�o��e#:+��E���| � ��JL�A�6�bs'�I�+DSkD�ta��Ο6��ܲWax �C��Pc�,�l�R'*��n���ć��B&���̮��1)�L�8�!C��J�0���މ��d�Xp1��A�[����͸�`|ͧF�+,}����@�za4�I4G�/�z�}P�/��^9Jo�x6Ƒ �J;?LF�h���s.w�	�f��s%/�%v��ٜ�]&Bn?t5���^�� ����_���虂ڏQ�/����>������uّ�>H���3���,%�"8H�A�f�@��2��h�9���/4�ض��P�:��@&�"��1�����yƐ1�}�r���!�������#"�1��ZQme0�s�_/��>_<3�����oU����On\���z�SDO��/ϱë��f	��ubݶ�Ȩs�MI�Y��머�����3b!�w�����x�B��u��O.����}�x�Y��R�%�t �-5d�[SH�,��X�W����}�M�Dqﲨ��G��H��
�����"$Ya��[�G6��ì�1	 �_�_t3-��wt�̤Yn͹����P{z�0�֯.nQ}��zV�$�D,rڹG�t�����ȾGf����F��#��c�E�3�1-������r9���
�E��ږY�P�w����J){侥`	D�(��C?	�ڳZ���
��4e���6d��@%�f�%���B�-#���Mky�Ӿ���6Y��"AAn�DhV����w�-����c���o���^Y�TyQe/�?%�&��O���׾9�#��[��EES�����B3Mzf͌\�[�C�s8op}fYE6�S,Cq��<�؞���Jx�����?�)��=viG v:�z{~�t����7BI�'�o���Xm����2{snh(���""ߍ������L;���@q<j��a�R�K��}��?�����>H+a����}��$�`��P��8��MD t��~���4��Dz�;��-���ۡyfO�O����)3��w)d�� lʧ@�m�s��U'�#K�qe�/�(��q&�|�ɱ��+n�~��c(�������9~��+fi���Nm�`0h�k2\������~b��EwD���G����sQ�.�y/N��S+u-��������L�{1�|���n��2�B�c��f�=����nT9�i��4p?�����<���i�aQ���:A��C��1�X\(y�"�P|0�(gͱ��#�@����z<�ph�W���Uƺ9�]d��p��Ȟ�U\V����l�ghms�Ѝ���mF�v��	��C��ߵ#�8�n3����5����u���� �zχ��ؤ��!]�UE�����r�E�-Z�O�5a���lZ(�:<�׬�,[�e�Y��ŧ4�84`��p����6��1Tչh�b���I�9��7+�@~o� ,���JW�r"XS��M�F�1?$#[<�� �4_�n�R2��Tr��VP�%q�W�f �^I�
Q��QΩO;����x`��LcJ���˟1JD�̐)����Uue�P�)y�/�o�1�lc���C�WO-�+�]rG�%�A �����V��
و���F�b�]7��������5��/�v�K�EXߞζK��m(�	(�z���)�� ��O<�j��*ޢ8L�-�5�,D�o�XUH��3�I��K���+�7-�ԯ�L��.��;RҨ]���oL���~%v@�T�5W�\�t�s����E+��4ˈ�F���t��%�]H&}E�ʬYIv�jG)CUBD�
�x�&��/�	s�/����j����[��65����������\[}I�_f>�wԺ�U:zZ3lH�彫�����j������������}���K�HP�#WI7=T���+��$z�8Q*o�V��Z��Հo�7w�"Ł[6Q���'��2��bZ����:|j�����(C���qf�>����MM�u����&9��pk[u���!'��7���ac����Mr�87��~��!�fA4BT�����z�s���.���cmT��!]�1�Q��T�
��n��t����Z�qoH�Y�����}sZQ�R�$��@��������s��7v���oS���04n?܍q�X*��l�2 �����z��q�#��kXP�OD;lY��I�����ޒ0�H�M�����LÔ�w��(E.;6AiK	#�hq8
hi�ԣ=�LQ�8�fBs~��3/��&D�8|��>i���Fg�R� �D�n�ۯ���U4�<��5u�~��,�]xIg?&.�Ud`��X2o3{�������r��_�pE��w+���� ��@���b���f��N���.:�!9�b�Q��a.fe/(s�ܾP�t���G�1	�cM��li��u��
��RnmBvrʄ�;w�����^t��k;�r9`zny��Cl;G�Z�i7b�lq':�ť�=ޙ%ц��f2�ϩ���7��/Ю�`���S}R�ge�W��k7�ѭ���͔55Y=��|�Sr���M>�^0z���NC�U!��_HE��k<:���2x����Y�M(D�j�̵C"Ѧq3ϊ�`�Q
\��,hZ�d�3�>p_9��x����ҋ �����^惊��.�u��=i�ͻ��z�C�n4 �{5�B�]�J�0Y���OU����,�����mVج>�:�eR��7s9�K�%h�����i��q1	&n����
Q�s>�k��$���5��e��O.-n��f*�*�7�d1�l2���oE3�N~��u��Վ���=���
U�|ٓ<��e���/�/.Jt������z�߁���9�
�5�.��y����JG�V3����1��}s�H� ɱ�R�T��H)_�B�3I/��y��A}�Q*�Y0�p�E��B��;��-�%M�O�������s0�g�g�-�Y���zv�?L_｝�J�R����RA�	k�AiK�=C�Y�����u)Q�jQQ{P�9��!|+�	{��Ǐڰg\	�~Q�dw�� >g�R�k3�-F�l��$�Q�V��(k�������%]XnI���p.8ɢc�D��)\��D�>�y��i*���+ar��X�'������_ţ�z�r�w# �\QS$���$�2ȁ㠻#ꤣ��~��Y[X9�|,#��5⵬��Ǘiv�tUt3>ğ�1��;98�05�.�#HcxT�0��?_�����̖���>ɫZ�ޓ�Ս�)�]RQ����]�â��Z!8=����b|P������}a�B>7Kk�2��������{�S����ľ'�X�a�O�<�U*�Dyb�X���*��5B������~h����(ql�1 ����s�鏏Km
�XEae�Ϯ�;�$��Sw�:	���}(m�<SF���@E��,	:m�+o���2aR�������W��G=��]\�1�
����s�������YU�W�n��i�è:�h�/�d>F5rʊN.aJ�04"���.hJ�-ώ���Dg��$�+���K
�s�Z���M�(�>�`Rd�z�Qx�w#ul��7\��}DލF�c>g���]@;Fq����]�%����DD"���ۊi2 ���a��1jW�G�����`e�!�/�Vr�I����ל7֒���ҝ��cNJ�Q��2D���[#J��#!���y|��L���ɡ�b]����k� o�]>�1gY��X�R���77� �Pa@� �� �����q ���e�Q� ��[��<Y&�Y�m���<�~v�Qͤ+�E��7�H��\�?���c�M[8�)	�8�Ѳ�$l���qT����P�h�������������,���<���~ҷb��߻ݐuh
���^+m���
@ȷ��|��S�5}�Ǌ���A>���e|�9#2�G&�|jdrz�OC
Rj�O=�tW
�̩/,�����H����$�P�I''��ީ�l�Sߣ>E���H��b�C��H��ͪ��[ǠR�������nB>��[{�b'B�sj0�ң�%��e\>>I�ß���ˈ���/o
y�:{4�jҫ�q'!�x�w�Z�M��<�`�!.R�����ƾ��D�V���D��2��5ñp�K�c��G/+�����ԣtox���Н����w	��E�q]���_i�®������-�q�낹��c����TTL3��0 �U�R�|�7���#+}�}o��6�zs�+!L�2>!Y������`��tT����3<ZI�I�~Zzi�e��}Xl���P�mH�V��T����MY�>�W�:�{'�ϒ5GY�a�F~|S�3�ڇک7آ��/�<��Y��l�������J�a�ʹEN�*H�����3�q �.���6�C�1��ޗ7is|ȧ�h�Wu�E���ǹ��S
R���ת,�5����J6��5V���^�"4�h�M��P� ����s$�3ΡR[�O N<)�d����
���8�wx8��8k�P--~���}E�������;�x~(���.�k�����Z���1ya��&�H�
��yW���ń�s�J�&�@ٖ��lf*P��if��̄��S��]]��yo�3ƀ�1�8 �V��1���E���s8�vg���J�Ŋ[�r�����̊_H���)#c�V@��&Z�>.��O�͓�;M��4��S���SRȆB%�@�`S�l;
#�i5�uސ�����=qٙ T ��=ȽK�Ԝ�	��z.�c�3� v����q9���\�c�g���=K�7ݏ3�$�5�H25~*��	�d�(йx�:`ct���j+)�J�(/7�vB��&$D�Y<�y�[NĄ�ٹ<��p�ZH��ޑm9����m�~�p=k"������!#[~���wF[Aػ	�pw��E@�b��i�;5���a�,]Ɍ�z f����j1o��G^{��/���P�<�n��ڢ8_��S�%{&��w���7,�]F*~R.a�'h�K��xJ3��ggW@18�iC1�f3���F�~�C��AE}t�ۣ2�v<�O$Ygk|d*v�X�H��0�MڤM���M���v]x���� ��7�y�֧��rep�j���e%�r!`g\qzY�"��?-u��6o&����vݸP�S�v ƺ/_�������]�6d�t@�\z�A��D���b�<�����Y� ��^������o��JzsO�h%��k�WjL��J� ��0�5҃ �����?g�!�������Q5r��~�b��f���)r��֡�;.���q߀�����̵+�aH�A�s�s��d�,0�תX.y䝖�Qm���a�>8� <�g�� q���DjE�A6B'δ�pd����-��܏��9b��C��C�M�e�f��OA�DDr�q��®� �X��)���Ts�_6wB3D$�O2�'AҞG[��H�9��*�ɑM�]�)I�;��5} T�*��qNqc����AL3�bu�d-D�<hԤ^�����3����7h�]ͬ��P�WTI�'ٯoT�K#��>(�f�?D�a�s�t|_k�n�t��_��HK=9LS�K7c\V�}#l���$jq�%j�@��p��[4	K��p������[�k�Uvn���?�ȷLm8���ZN�W�D�9i��o����6��$&��a	PP2N���#^���q�ыhEm���pZ�ʯ,�����	~�Cz�����N����=!�8�8;7��2fH��2��5(�[�Ax�`�i�c�dg��͌n��z}K� <)�@�Ͷ��^n�)�߻�i���/keW,j~<���UF���U�%�E������U%KtIg�.�栊3n8�ɛ2������_�֣~1P�V�Q&ݻH�S&��04�y+��p�����J\5��
��1��B����3OA���]iYq�V��P�m�3^�w؛���Aq<%P���.K�\�M=�{ų�l����D��Z�h�B��B����Lu4�jzY3N�s��Ú&{��b0&:��<�������5��������Q��"���K�������O��t��Q�C�Tҽ��QςHcϥ�#�N���cцqV���'���6�F�Rb�_��2Ir&�bX�1o�ڜY������
+���;O��H>I��N+;�a���[#�#�KE�x��d�Ζ�1
CY�pvE|�%��I/�O��XWKh�i+;S"?�e��[�'�p%V�pI�ȥV�� ~�(�_�F�|ru�ý4
�9���q���Ågu��b�SLm��#������ę;%Zb�x��h	E]�f��j�����k�jo�e䦎h��%�O�}"�XH@:�q�A˃�GC3�Ia��=}��p
0��!-��z:΅��^_�b!�F��wý�Ǉ*���m(h�|Q��u�R�"��\�R)�N�J��w�����Q4?��Mh`���:7B��S�`��i� �mH0$��?u��K���j��4#�%ڋ6�]u|��&�cm���\�./p̬"����y�)"	~����"��{�f�;^�6�zJE8���(�d?���W����������U�,���3@�8�&�K�Q�N��Y�qT���߄=o��%���W3$k��,W���^�k��� K�}�]���$�_�l�Ê��o.�����I�1�!`��@{bme�����Y5<5�ܪOB|��e*� ���9�L.�I��%�[g��lv�ꄞ��.,�K�5�j�N*��m����cԄ��뽗�じ�1�<����f���0Z��W��p�SND�Rn??�o�e���8�b��6�
*v$p0�}N'gs������������)%1�0�sؙ������8f�q�nP暷 �#��åt����!��f��4x�ʍ˧�ʰ^>��ғ�	��0�f�S��h{�}�C6�~��OhS�p���[/�;ǘ����ǟ��u����Z�[��G�8��2|�g��*R�K��ѽ�Y ����L�JƺF<Nk�(@�_�o�E)��%Yc��L:Њg>I�IMmg@Jq�)]w��8ޓdĢ*���%�����ZS���x�FT�p�)J�fi���K��b�>�= ��"/`���l(g���p#\���⬄UQӧ41"�ڍ=��gu4�P.�3 ���y���ɭ��Ւ�=��0��֜_~x�T����R�XB��*\_~}:��|D:V�F�eF�E�Q�q ��;�g�2��}��9)���1�����)�-��Md�S���A�
�|6�lO}&%�ٚ�P���������&$e�
�W�D�ӷu�;��b���}L2��S��&�4��t�9�Bo<C��ɨrϓ���XIR��ˌ�I-¥:����!n@� F]-;�'Fv��7�Qr]�������3 xtxo��M����P��
'*��}�i��C+fZ��Q(AA�!~M�~X�^%�1�AC�r`}RT<F%�Y�YG���'U�GQ��}/� v#�*��ޗ�^���u�	��( ^�^��צ���^���WZ��ؾh���s�9�W�-[��g�d��x ��&f���X���QՒU-�G�v�'l������v���a��MT
��d\��F��Dʽ�a0f�U�NV�
�-������e
�Q6����_s����u���\�[X#���\i�p�䔶K\�q9,����\���3/NW�]��J}��C��Wˉ��'�M��=�HV���?#�1��A��KJg"�:}x��K%�`N��(-���������8�����V�:�|
�L�=��NJA5�ڤڹŀJ;�5���2̷ �)��1��?�̷�D��E8-�mt��è�͖�&�uX�qL�HL��Zѱ��\yb�@"���saP68�^�u%E�B*o=�K>���D�<�PoY;jKC�J���f:�5�jxT��!gޖ�HG�n\��y�:�d��5q�͛��k�6����8�٫��0'R+��7��$3&g��8�*�lw^�����(ǣC�.yq�
�����������Q����T)�4�%Χ9 gz'�����Q�{�-�x.s;�&)bXK���X���4��}.#�HT�H�S`�	�F����Hu)-���`�yA���H�@�[ۓ�����	+���&S�Gg��n�-y�eS���1*��4�������d�"J��5܃��N�m�	��o�E�r\�=kV�+.%A%�祵�!�@�~Y���j�2�(����;A��P���t����f��z��(c�ٯ�q��Mڥ���7�g�X�#�Y�����o���6�ޟ��\Ɣ&&��"�oR�m%v�:v+a(_��ؤ�ӹ_���Lٮpt?AH�����f�Ȉ�����Cr�@)D�5�u���N��`�ЖV�;��#���1L��S�Xj�9���E/���7�z���oj`C!g���H��$�.�E��&� ��>�΃e�?i���W�g����ӗ�_J�[r�*Ĵ����B8A����%m�AJ�����\�H_�S�,��</eγpJ���U4Eޙ�\�!��T��k��Ȫ}�����Odm���W7ӻe41P�~i��_Q}3���E^l�n)��I1�ʹ�r�Nٟ��.1 �{U3yR�5��hk�5�7�+h��PV���6�{�~�o��g��+��#��7C�@]&i���V\����{y[�>�N�`�h�� <��K��}3�+��c����"��� ��u*0� _H=м�&���H�m�r3i��x��?����s�S�߿F�ۀ8{S��a��(zidbQ���xG��[�'�O|�@�z���WsBW#�*�t�@F��Ѐ8em��{j�m�003���I,}ݸd�e�k����x�2�gt�쐃x_Z.�Y!��N�H�B�ɯ�f��י������.� �P���5̺��RY�w^oJ߅�!�~5Y����S��9��!(�@-�s�lΎu��϶�vg�ޝ��v˻r�d�� �Ѩ��$ o�8}�C�@S;�te�,�c4{|�s Qb�i�`��f�)�F��F�/!�=h�bƜ�q��0�l�{�pS�)�<W�w�X�D>��@nQ�-t��%%�� 	rMs�w.�JޜH_��x��hߍ��G��+Uϧ?�(�ʳ}��ͳ|�};�ғ������Ͽ�^.[z��� G���������B�"B��sډ�S~P��$:[��:�� 
�yH�D��|k]E/Ń��rS�t]:�Ѱ�K
JH���Y�`�$|��w��J�(G�ʃ��+����8\;;��oNRh����=�(���<z6�:���	ἐnA`�#��W�oI���t�$����2AXZ�E V����H�E�Ĵ����0�<c�_�H�m���(�`�e�&p�P!vx����3[GݗtO�iam�x�Ƥ��Ǝ�r����h�<���ǠrFwK��l�=��{k�~�X~q��~=E��|ٔ��k*K?(;�D!��ղ[�Q~͈Ǒ�uz[�;6�⏶�3C�u�]8A+�Q����ᙙ�I�������ע]�E �P���~H���`��BY�3�H���`��³��3����\wL�fA�}��գ��6=�R'r%� �E��d!VYc����K�>E�//Gh�[
�<W���!4΁��~S������:�Fo�5�����f&�v7�e{�H*������Щ����s%F�B|�Dk^��e$�d�ja$ƦL��,_{a��К�&�I����2��V�z����������ɟ?����!P׸{]��spTnTf�[�)M���K�p�Q�@������2A�(�
�	N��3���a��`{�̭�H�Oyd���|}h�麟��0ljQi���4�{E��z�Q=��ژ�[#��O���!�O�r�[��C�{G��н�f"������d��7���~
�P�����>4Y;Sp��$	���R<� Ae(#1yBjtR�[`�a�����U��$|u- ����*CN�]9�p�"+�~�^:�BYh�~"�.��7���0W��e��QJx��`R�l���,B��7!^�c�.�i�e��T�U���3[}8�ĸХSs����}BKeO\�[�sܮ��Y%*\�;<�C+��/ڋ���I.SDo&T��C=o#b��u���k�5�uw��B=.
U�D���Xz
��/e1�z�u�y�d%�m�V�i�B�S�B��z��������z�qrEk���˪�z�A8f=f��n�q&d�Z�F�D`��u���U
��tzP��g��[~V2����X>�L��e�+M��Q1{������:��!w�E��kv+�#��@^�ܪ�Wl������/�^1��b-���N��w�)��:c�~�\'n����J�������Q_�2�I�ڀ_�sw���L�z_�����,�tE��n U�u���0�~�C��')$ʼ�y�4eݙ+��<�K%��%� J��z�磔v���2�ܳ�Rż��7��g�q� ��$�1�Icw %�������������c�o-��,��f�s�ڠ3�PV���'��}�WPE�
;D�4��E����D�p;�Ç-W)A��7��[�?Kw�j��D{����ѫ�r���X=GP��1�m|�.W		T%h�Z7N*��h�[F��3��`���A3���ǰ��rq"�Cq�`�?�ؠP8��_��"�ɜ@��+���c7�G�vo�.sv�$��� (�+5���y�5���s<cpk!s]E]-�xq�h-tݪ��H�(N#7�S,����I�H��e%���Y:���?�k?s��Y�%K�<���@.�q4i���8�j6�>U��>�xA�8��I��!��X�x!��Q
���]bp�!qb��Oݜ�-"����NaIޞtrl�DČ���ZF�&�ֺΆ� �T�����P>����R���S/P��̀�Y�և����,˷lEmhu�������e�I���I�>�w5Q�[=�Dg:��ix���Dƛl�.kt��r�P��UAbۤHF�����ZF�����l����'��@+�6G�:��T1�JaQWEX9%'�|	��m_�}��Z���y9��Θ7���s:&*����XH�d�//��+G� -݈��ű�>ɨ����q�qz��1W-�Xx�jt]XqDڥ5�O�Q������˘�RG�& e��3�:�8�ʒ�PQ�P]{F���R�O�M]��\*;���[DN���љm�~�!���g}���T��p�5���?���$m8������a��%��V���9���g��t�t8a(�[����:L��C�\\�*�6X�Ǖހ	�>h�ߕ}K�w��pW��ܳ��vPRJVC�yvg�{�G�F>͠��8WW�(����→����;��צo �?�1�
�ڭ[��dH�M�9�hl�� [�(��{��<}�O���H��/v#��U�M��R�6u������/�I���Co,�;�^�7�'���9�[3��O;o�M��
�2rz��X0��t�f���t@b��a��3���n�76�o�I��;���Nd�m�!z��W�U��T�������=�����,��T<�ԅ����FP>���7��R_��u��9ڰ_"|n4UT*�@�̀��<�"-��|x<]�U��-���u�TF-f:�u�0QY� �*����4!c�[�<��~��,9�w�Y�6����'�<��I��ejwij�~M��)�uu?�=���2d�)�L�1j��w�B���� AEu��u6}�OF��F�����bs��͢����Q/�m��<	�!�6��u�� a�/αG;�\ƞK�P�A���h<�AOc�x�Y�{>�:��%��<�f�e��э��	һB�'��he�K��yM�븈捄�3��|�M����H9�����J�HC���W�"��b�4�Yޒ�i��&&�LC�Z���%��%`�b)��^����W��-�?޿z�,藰� +�T�가qEՖt�x�i��x�Ր�Z�lΩ�hx�%�[��b�v VRVKnD;��c���ڥ�L�6i\y2���P�E� tP,�)|��-�<-_1
<���GS6Y5M'`���p��E�9ʛT�q��.���QZ�Sx&��3KD��������c�>Į���o�y�d� �w�3�`�Jy$d֊�Υ�@�ɪ�����ԿWpA�Z&��?�9�Sww��@BOD^h�N�JQ��f"r�Uq��c~�
��
���S��:�=�P�oW^ "?^4#��Y�D����)B[��s�;�3J1�n��������)MI�,��h/�{�P�j)�/n�@yI|���~�=(������q9���|?�l���q�@�"7@v��A�#!+M��
�2�K����&�r@X�.�*��IVkyH�T^A��$Q(� ���ֲ����㴙_��@�f��.U�j���\���;��$����`�,��8'���1�� @x�l�ʚgO���2KR�'NL��Ev[���<�@�sA��|�}�A�N���)_��Hc��R���a�I)�Y�a��g*�-�"��y`_N���A0{%S'^qN���&����:�z���l-�W�ҕ'���< ݄��؂�aCH�o+*��N:z�f��y4��&�?W ��w�,����<.T�_�	�z�5�w,�½윘y���uD�mu��82�u2�W��������	ύI���f�-c�?�4����QYA1އ��\���� q���~� ֋U��ĒO�j�[�q�������
,�_4MMޡ�d
M�{���F߰h���h1�����o�RD����Ω��p�g�k�&�/"d�_x����rl0 �����PĻ�pf!�(U'~�Z�£���vƓ��=ܞ�o�,�-|��g�D����|lĐu]��O��>D�C|}s�7&�<�W�F��^
'��M"=W��>{J���)���L�OO�f"�E�� ֖Mb;�0q��,�7�c���P��V *z�1��#��d���ڗ�S��OՐ,3�e.���`{M�~:�79�K�δ�f��mT�%�fD�R\��^?�`��n6Kz�Q�r"]���D��S,$�vNs���N ����n�V��ȣ3HD���ȃFi�i��X/s�.m�K�������.8Jd�(`��'=�;<�i!g's�R��b���P�K/���-�S�k	[��p��&�����Yx�:��}����#t	p�]�s;�^~ bp�Cw�Z�y�?�Wk�؆,ĒyeM5)����WG�[�1���Z�d���v��"�ˁ�����=�Y�ޓ��	����m�1��i��ل`���]ǙG�
&B�MX�2���@;!�u�T�Ѽ�N��`�N�A�ro��:7��b�[*81��E����+{މ�L����++'/��^�>Ez}H?� WH��HED	@�nx��1�#��J$x�Q�����wuHA�!A}��p��ؐ�͖�r��I�Ꝩ˪E�,�1�H{��fA�lPX6���
,�ۖ��ԏ��p��z�ړ�?ˈh��˒(����c6��	�J�:�o�9���j%�QzBL=�֦��]q�ԍbH��
��1�`�"�k�rc���F�'�dV^�T��G�m�un��� H��f��1��h�V[k�t�@�e	�0����\��H��;_΁�NW-��nmy���c�f�<��`����AL���@ܵ} Y�� Ϝ.qBC0�0�H�$=Gc�c�����Z�~hay�>���vUU:! pM %��x/~�G�|�I5�[wV�_�`��f���[�Hg���n��&�ێ���q>,��9�����1O
,�����᠋Mh��i11`���<@��@�>r�a7�l��/ִ#'4�Ě�}P�=J���w0����?�:r0H!���b-�����-ٖK��kr�ē��;~<��B][�j6x�f�cYA{F�u��g#�PѥD�#��F�
�;����,�\�C�:2�KɽK���v�ڗe�M��(1n�!�e�8+$u #�u��я{��Lq�.�[��~���-�~2��x�K ;�Z4q��uw�<+���u���Ѡek���.ٺ�˓�]��_ X��K�� ;ʧ�l�v@�[A�:����Qi�X1����}ͽ~z)���I|���|I0�51�@5�#Q��ԛ�vZw�3b�pJ<��ۉ���Ox!<�{m5�1p�8��f��߭kd��e=�CglE���w+x[��6�*�]��y�U�XmQ([�Kʑ��nT�5�������X�v��ͅV��Ѐ���Y8yS씍��� ����P�@"]�"e��mKG�]�2�0\�CI}�@�[kO�Ʉ�|[ן̧!�=����Ex�y��d����ٶ�+���6���|\���`&������ݺ#�q�d�6�!��M�LGp�It5<�W>�,��&�zbb�ݓ���o���	~�d�,;�:8�H{[�-��7�0����k7�U&�N Y���|kT7�(�=@�Vi�/���܋��CXg}A+n�dy0���g4��R�:�mU�bq�h�#=��M�;��#�1�!��>�;�R"���t��y�v+�B7ҵڞ�]�>Y�=�v���Wԧ._H���vn�w��z���9�c:��ԗ��^��&�ׇ$���˶�*�Uc'��`G�#�=�8|�+��ꃎY��8�*D�I�@����e=����=����`sK|�tě #�))���L�V���qת��n	̍y���
�����$I��*�%
�f\�D��X_�>�K�R�Y^d�<�%<�%���B���{�`������K�#?���h��y�9�K�6�y~�ܠ�r"6e��]�~���Ew�R=v�7>���pZ:�j��n��~,�6���4&3�	
P�U�'	��]Ui���v'������Ȣ��uU�/_H0b�a�0�������<AKԓKڜ=���|V�Te��,U'�n�]���J��]vk�-F���TC?��s��$!���Cƛ���W��A'�z�0tS�ϯ�JB��Z��"�W~8��*��QU�ԫ�l�X�&�&��hbn���*S�^�
�D�贺"�"3X��(O��3-uz1��Ϻ}���)}�b���zսj]�s�8�Y��p��k���k���j`�Y{+l�a�È2F������Z��a��ϧm�.���������[m]��C(9N�r�S�	j���^̬�}���r�vrY�t0��V�|SW����S�J�EgVa�qc�q��7?i���pf*�NGl������Nw���"��'��c�,�aN���6O�իr��B��+;U)�ѧ8��[1�DW|xĕ?$���ȃ�+�:$�#A.�u�Ŏ�J/#����3_B�ը���X�cN/���y<םG扆;�Р����FV�gϻ���A;�@3��1>V�T������Cl
QR�N�_?���e=�'�q?v�0��ǒĄ��؈����2�C���M�5��u_��{wiI�Wz��3�� ᚐ��g�!
�*�4���Q�ևFt���ݱ���&W�x,������)�f�wm@�3�kFyK�2\j�=�N� i���/X!�Lm��[�JBU��I��3; ]���	
B���	�6����w{��{sA�m�ыm�W��%	�}H��[[��ځ��
�I=���t�%�͝�'�V��!��|�a5~;����O�F��es��sǟ��X��t��7B�G	w\l�|�N�����}������"�;��kI;$�+/;מ �ʴ�L�G��l��i�~v�p����o�R���F�2\�-�4���}�o�b�*��,��#ϊ&5ԍ/��;]������Ӻ��[q�0�zG��*�-a�Q��#���|7)��R^f��}��4J��@n{|{��@?ܝ�Ӥ��)/P����Ҧ���M��������ڔ��{�r�]�]��a��K�6�i����I�- �<l�s5@�K_���8,Enn�LdG �;m^W�W8G�@Q�q�4p�$�x�q��r���j��7��ˠB2�wgf��4;�����ñ#Xq����M�A�yf��q�mB�������_�m�M�vS�jIUC'e�m���=�h?�e]��G|�����Q�9w%�+LWET���E�@o��,!d��JO�;�s"v��K���3-P����)2�@)�m�+��}.Y�x`"��6c2%l	�,�)����8캋��9���nfT3�� 7�;�E��R�(M����͸�����_��:��6
�s`�(���7A�ґ��Y�xԨ����� A9���B�e�jeB�d��.��|k�_�H�a4C<���*�|���m�>H�P��.��Nk ����j_/�k�H.bU�<���M���л2��S�ާn�����-��L�i�Z�>_���������'&��+����Z�"o�2n��cί`c��[�
����(9�vm���{c3M�����4K�R�G�	�u��0ў�1�����p�e	��$��T�Ӛu��O4(e�#�}�#ԃ8o�{��6�9,��& ��P��-�ދV�|^2���,M�e�Z��KT���S�nM��"�q�� 6o��>����Q��M!�d�k����	�^��cf�[����@q$T�zb�,������l� �/<����.%@��h�RH8#��զ���Q��0���?���M(��.rSz���[֍��~�8��=�<�VH�����'"��zc�u�~ø��#c!�	�D�y�/�����G /\�$0v� ;��cQ��:�t��	��`B���{'c��YRcom��*v��n�����1+!��e�&�n�!���)5�(�m�p+t���Z���/�X���k�Sr a��x���y3����.N��J�æ�qR������`oՐEF��ٓ#W�"-3�w�f����D�lJ�d��&�_g�i�Er|�"&	��(���(+j:��S ��`�O@J;zɓ%��f>��tg��M�1�<��6�]����?/:��]�3�PD�`K��ܦr7���8hb��+O]FZ�-�j��Jٰh�x�b�pM�'��(�^��n����@ZVz�I[t��.5�;�̎����֔�o$�\do������l���k$��__��sї�U���.Ҽ#��@g�3�\Kɲr�t��vz5c"��q\�է��֖�S(�K�P^]��!�p���T'ߍ������е}�@�)="�w�5���{��_�}�·|ȱ	� ����;Ѷlֵ���J�K�o���$�J�Wv�Eן���Yl�!��!��-���q�NH-��+�tqGy\,K]:�
��<#��X>]�S��v���?ÂE|K��gY�1��Ͻ�-M_]��0�)'�Gޥ��u�"H;��8)5�z�(y
�X@.(���ux�#�S��A:�2T��ћ����(�d�w���������rيD�[��m�G~/a��Ӝ�WP��mp�
�u�`����.�]��/��7�/��d:��pL/�[^?��ƽp�AAAh��+,�:��O��g��Lqn�x2�����df,ɯ�����,��ı�BCfد���vg�^s�� �E���"|�U��ڽ�)�@��ZQ���`�L/B6?H_�V����ʣŋ��2,-R���.b}"��[�.���۹�N�qGe[N;�/��a�l*�%����y�uPD��
�Q�1*�`IY��K��mj5x]����V�#���/��j%"�����,��Rq.�0�w��O��q��';X�e�����(��G=��ب�Y�{@�I�V�^l��b�;�4��.,�ƞ���E�a:�&87`!��*o�m�P���]�t���_:?�2+=���hv~-���m�?Y���'��(�,%�z/����W}�$���ǁ���8DEz�>�3;,ܾ��I�I��b�S8c�1w��=>���[�2�.�)9�~]��n�' �x왋�t�l��g�Chu��FI�N<�O�x�c^�
�C$!��V�^���Xث料���va�,|� ��(���p�W�m0X��nY�Fy�ȗJ��\*ax�f�W�f"���-��H��aH�,��j� Vw�%�|�A]��=���@�cZ�ҭީ��&V������M�u;�Ǉ���@8�o5�rT,.]�w$-cc�c9	����J���'i�?��.C4�l�R�n-��ę��cj�%J+X���:N"2�����/��
,�
9)�I�l�;ae̲EM�뉑�֤I�)@��]�1}�Zr��v+�A�4�b�ɡ-m�	]+�M�<3`����y���U���cr��t	�= �陎u���OX�؜�	M�*NN�)����7]B+�G���89��X��G�U�;����1�DL��V�CM 0d6�d�V7%!T����+^���n�H3���ֱ�����$/4v
�����g�cll���jvI��A�3����@HuM���&ϔ��Ɨ��v9�^G�e�L\���v�����Ɍ{q��'��>��劂vBţ����,�"M�9y�l;�h��4{��H)�6C=ޔ���L/ܞn
�n<�@3�5��v��R��� y강q8�>�W����X_���:\�|nb�w}p:Oa��Gv�)��_�d\R��۫��T�"0�
�#x�7Mj��_~�7��ɳ�*v�Ӟ�;"�����H6s�m�W���%d[6�rx`H�^�*"��૝YҖ[�Ɖ�D��GƏ�����k}v�0���9,�#�G�qG��P����|����a�?����H�j��W�	P�<+Ek(mB������� cͳCW��8��e���7���G;��?�-������%�d�� Uи�G5W��=74oi7C"�&�'�Ek��p��<�m�[v!bG6�(�,7�'�Y���ڮ��Kh���ZV��pp�-p}��!3j��$"̏�nO�t��}h{W�H���ْW��QdJ2���ynpP�:��~C�ܚ�@;�`��
/�2G���J��{��d�`��d��&`V͕0ъ��+�עt����	w��ͺk�X�}�7ݝwʹ�3'��J��*
r֫�5w��R���N�
ds]q��J'1l�1��e`�j{�ɘ�7�t���kf��pS�3{��)�]��NL(lI���3DӒ�?�a�>u��}�� Z�hk���lz<6p��e���	G���6ԑ�ө���%N��/ �����W-8�k�F�0��(�{:խ��'�M����@�4y(?e�^|�5���F8����W\�V1W�l֕S�
s	6������0� a�1Dn�!���P7���5��"������`��@�o��j�)�{5���?����?��N��_p�c�}����#\n	xmgʄ�ܪt%%�\��b�l�\_i��-�5A�G�Ә[;�gԮ��ε�VY�*��E�]X�K�Iz�;bi.��%iפ��p"Z���G�i !=-N�E��`��a�7�4�S���D����៯��U��\{x�d_o7/��PS,�K��s��,��}�貣5��P8���f�JU��Kޔw�D_1�D��k�_7|l�2��N�G"��}23���Z�8$���s8�L͙ԩ�Ls�H&�!*MXD�D��'����6�w�3�u�$^=�p���99���8�R8RM�7}x�b���L������+������x)j)D��,�!����ב�(�٩�v���O����!���g01MZ0F��h��R�"_P���ӑq��&���g�G&:.k"�{o8K� �|���>��/1dC!���l b,X��u\TI	���pz�U��8.Fm?CU1�F�x-���C��.��Óx�u	ܦo�A^ߘf�am�}v���3dσ�Mxw¹�>����s��(�m�Y%~�H'9y�,��v�^������wl O��o�g���!2;ᎹA$�,�%H���b�}�7����H���/�(ѝ�2�rx�˚�4�,{�m�U���@��R��c���O��HN-�$O`����J�T�'m�	�wf&2o��0"~\����I	���7�+��R@���.���I���� y]���=���KUCo~�`*,Z0p ����ɆP��.Z�':����5(�f�+��x��[!E�B��.��y[�d�(g�]�|Ѷ��*���p���@ϙ�N�.#�BO�L�.%h�$o���8���WNn8���Ud;5rA�
d=���XfXi8nA�Rx���1���\l��|�$�)�z�i�W���Չ�|akc^�v�3��6$5"���*q�l;@����z��
�um����p3�١�>���fɇ.��
BN)0�<�vp�I�����1|����|Fd���� x9�x9xoN{OI�Z*��
J�}��݄(�?�MFE��h��<�
<�������7Dh�3!�=�;�F� b(d�N��C��'��U�b�.)����r�6�q����Rt|xIZ*c��^Z��fqˢ*Z��q� :������*yM�΢F'��H�ټ�~�Utg_mFu~��<�������]��뛰�k����	���ZS�wV/�_��ϴTG�
�|5��.�'���D�8l�ddF��Ω��Crv+y����P��-���4!���2�S�VG��"&�.��(tTlB��/�	�
�jTM&���%����ȞȀ��V������y�����zO�)�� �����������%:Q�����'�;l�\�� �z�d{���J;<�WqΩ,�1-2S�I�V�%̛�Y�hd��X��_�ڰS+�iւ�����ɪ�;�*ܙ|�F�	΄d1蕉%:��O��=c�`���3�-�B�LGh�M1����N�A�����^Zg���ص-;rA��Mf�-�L7��KVIX�K	%�<�w.�f�(�ۈ	|{0�����>�t�+����`�q锽��]p[�-��ap�fО2����y}/a]dK}���5��[�D��kBU��9��� ��j��:��~����',IE^n�F�C*�Գ�>M:g�0�Z��ݸ#�%�^�X���?��1�R���(�۽��(��0i@5< ��ŘFEK$�=��F����4���ū�|���!�iɺ� DAo��ف�]\N����n;��'�C WO:VޓRu��}S�����xc�QT�$X�i�W���Q}s�c�pF/c*[G�w�O���I���V��;?NO����S��JS�@���tdT�W�|��$arV���7$N��8 �5>40���P5q�O�`��5*y#�)�ڝ�n3�bA���d ݙ���L�m�:}Gj����v�Pb�77㊮H�T]�f�ۿ{>��+TI���6��&MH
)2�B���Qr�n�1�L�l�q����ނϊ F��%�q��&�ig(}�0��t�zC����I�0dccųm����9˰$^8R�������di���� #N���M����Q�Z���俕�=�\�|��\Џ���O*~t��;��	��B���R�y�����&������ኳ��/�ћ���9"�uAC�U�j����-���A/7P}�(�?��f�tO���ݙu�Bi��x/v��+�yP�0u��i=Ծ{�(����ɯ�5x_�Q��v�����ׁP�a�+��#c2�1��T>K��ͥ{hO���Zp'��d���r�k o�cW^v�u}
vs��M�9�W.^�Ҙ���7�.V�<���ƮPgА� c;��[f�tm@�aD�[���"}����"�3e�g��ځ�ₓ�x{�f�(]A�?��C0�Nt$��26���Ǧ�K4��Is��)�A΃�Gn�vq��0S��ؓ�`EI��Z��yLR*�w^��h��ֈ�q{ �3��[��Ga��L���2�ݩ�q���;��?��Atm3 a���Į�C�-��C%P�Ӷ����h�3�V�~����[>����S@Q����I2�l����� t޴6�<���z>��~��@��|؃E�z�I���R=j��?DD�3͓֑�O��n����(�\^���/6��d���{AM�E�)D?��K��+��U��%f�U�|���:�<����Q�0-���R��2���h��P;���+�L�gr�Eըt�g�����Q���@�ʯ�:�:��o��̀���/8�7CP����k��>~[*�p�8*b[ȼ���պm�ty��Ws����P9 ��,C��5��E�,�{$ݩ��?w�l�l=��]ӝ�dZ�`%�N��oyadzM���@	�w�mֶ��(bK�3��� �v��|0���C�n1�����nex�
�� �V��0��-�g�H3�E�K}`d���F��b�� ��-W�(<!ų��xhlu��ط�����H��0LEg{M�-cmֳ�Y�R�&~|-�
o/��PlEA��kN�'G9��sPb��PV�"������/�]����	$�֟��1lb�ȫ�I�m����$dh&����(9k}����r]��+�̇��EX^c�w&�O��c�p�^��F����:<�vpy̮*��09^WmV� �k���_�-Q��_i���C*x�X ��cag�W4&0�*�6_/�"C��E�ŎR7p�Y(h4�yP���~da#]St˭���<D%�3�=����>�5�eU�&l"�L��k���)�!�V[X�Q���`�n%����X��X(�,�W�c�����
�I�֌wA�q|�p�7�S�A�����R�q��`D5�]�6ݼhB`�Iu �$5�tI��,N��(ljWusNʱ�R��<1��L��"��kV��S0��-0f4��q��m7c���d[|�!�һJI1_�HƑ{9��*�p�/�1(~�����8Q�W�l�� �F����f��%�i���ߥ 	'e�"���?t���rnhҤ�
>l�����+<��ٗ��+<�l��j�"�Qw��3F{�*V�I�p7w�m�z&�'����%��Ѳ��<�a>$?��v����e��=��Ó����'�Ý�zw66 ]1�S� ^Ni#!N.q1���#3u�D�F*@��~p������)P�"Ub9�;8?��MO]�j����hX�P�v��-?�&��Ԯ�)d��j	�������ym��r��h&j��i��[�z��Dt��O��$��3�F@��w""��Qq�+f�]�т�rU����\lϭ�F�	�����$j`A�m���rxj�H!�O�q5��P��8�>*�k���;����O\@c�o��Qc$�Vr����?]��0�d{l�C��!�'�@�x���Zj��{�u)�	3%D�}��P��br��;/���L��"�_G�_dU��}����e&������q�t�y<�W�x�0����_#FNO�W��_ �?��_�\�) 1��TƁ�@���MM�����Úo��_R�VᵇEi_�0_�%0���u�.-m������v���R���#3qWr�ԶQ�x��9��B�Lq�i���#�&,���Vh��42�/(M��%�U"�,�M�v�������a'�4ȣ6�7����I#�h�=�z;2�k���X�%��?�����ve6Ϫ��t����R��0������٠u?��?+IM�	8��	���r3�}���e�v ��ѐ�N�1�[5�2w�
]}��nD��q��L�)���Yӿ��<�56h¬�	ԝ��v������H:��:�V�;��z�3��x�LWu5:�C4���m�U��%�=u\�WDJ�o�����2�B��A�3n7jeW�3���d�Na��x�G(���IK��4���Z:=D�W��R��x���i<�^���:	�����$mQ��=� D�L)� &�ʵ����F���Ar�|��s*�'8�˒-�d���1;*�c���}�f�Q�AC�'}���}�*��"�F��,��MkD�o�;�Q�,E2{�x�^B<x;}�x�@F�ϧ��ZhNĥa6�Y@���`�.��K�z�&f*��cg�O�l��@[�����ezt�N��7J���m�ƬќC�R'�����>��r(���ɐx��_� �Tg�2���p1�rM�b,/p�����^+�N2�hÔ�6��A���L�7s�нQ&r�"�r�s6���i{�SdX�M�5޴��\��������}۱Q����{F3�0�@"_+R��fI��X f������_�s�ǅ>���hgQ��>s�Cq4�:j�gMΉ�^�����2p���¶ˉYy.�H)��5E�No&���o��$x<`&�ݍ�Xc��Q N��<�.K'�)�>X�'�������C�VJeR�U��*��tr{����i[�`s��x�{�g�G)c�D"qL/>"y#4%�wB�W�b�nR#���b�P4p�Yb<���qp�}�Z��s���������4v�q�%j�I��'Z��d=��Vq@�8�_�����QG�`F_N����l!��B֌�cq�RpeF��=�q��@�8�����-��S�X�(���d�3��
w*f"�z
�y
e#��£�-�;}�W����s�ZrG��ܧ��:�^�u�7ɼ	_Ϣ�]-���#�z�J��rp�(#��rWHIO<IP�+�tY�G_�Z���8����(&e�������y$NY(2U�^�3��_�2�d�a��E� Ā2^a?n����:W#<ce3��+`K�<��J?�W����bJ໖B�]����>ja�#%*�=���H*��[���V�6>j��Wj�.!fܿ\؆����h�U�b�cyUt��C[����_�S׬GY)����!��4
���2!�E^Bh�@�S���LB��u�i@�c,��%��U�Y�AzB���ɘ�+]�z��.�|�%b	�S��;��{��3�F�h;���7f@��Br�poю����C����~���λn����zX�淚��0�Bʾ�jw��I�̊4����H,�NM�A������D;4�Y������
��|l�>����gn>�cM�S�����E��j/�N������>��lഘ k��؊�:�Us�{g��78|�?x�Oh�cڢ��#I��}��)��P�A?��� SV��G��%�g�8�� #/�ǻ�� 
�Bd.���Oq
)�\Z�5t���vh�lˮ�w6�d>�ō|�����CY�rg���$(�����on�|����p�X���=���P:2`v)�������օ�2���^c�a?��E�03�%�����~����R�z6��Pa?ozR/0~A�v�'�.����
����d�{x	��'������9׬���.�_;�L<�4Ό�6߱2��{0��"�c�ߢ1aH�Ƒ�(���j��	{�!!O�u�g	n�A�~�x]2���x��G�����K9ò����x!/�]*��o���"��Һ��g	� �A�|)eN��5 �1�b�K]�y$yk;t�g��R���úxp�A�n{9�H�~�(���[�p�4f8֠�h�dP���ᕕ�G�?Ղ۔��8ؿ6`������
�J��Osr	����$��Һi���;$y��o����? K������j����ЂLHu��Q�ˮ�p~���صy2&�#1�:��a�;�Qy�)[@Ny��2q�-O
t���4��k�FYn��f��5��jd�XY����bn��2L6�1т~�e$�����[E�O���L�1ǫ\��Ќ��d�aR��QN��3�rb�1o�.柪�O���1�a�=���M�h���]ߑtE�5�Mto��YS�՝I�Cy�˚��-���
D�I��)������5�oE]���u p��q�1����^ C�	�?�_Q-�|jܯ���M�?��G�-3&���JK ݿ]+O�����7���-p�����٬4�n��7oN�s��Ry�A�SJ5a�St ��2.�S�>+�O ��O{�p�e�R�\�J;D<��6�D(��w��W���@�a����yK��4ZG�F}�:ZK,�)�p4�ݾ�goH)�K��K���j�X	Ţ����xD��8�Gd?}��7����OH.�C�#7٠f��\P�1;9�����D��8���Jv/��k@gZ_�3��J��`.�|�y��n�E��E.ӓ냠&��7[B^�ҭ����������M)5��R�%a��H� �>�������_JD��{��ɠ��߼�
,���*�1lɚ�U`�Ε;�(�	���M�^���~E��E��U �U�M�#�E����zFFHu��F݂��jB����b��R�Ȇ���	���گ�e�'�4���Yu--���w҃�� 
CA���;�ęH��-l�������k ]��B��["$Vc�:�w�r�����^�8�R˯_vN�����#��̾��MH���]Zk��'��e��c��\R�0����^q�Y殀:�?bl�q^������V�W�k%}.���`!���G���dy1���/���2p����(EԲg5:@��z{�S���ܡ6o+i��V3�.v!ya�s�U8J�R�u��b�/�^����8=g�h!#j�t�!��]zd�ygor+LY0.Y%*7��p��v�Tq���Vx����.�GLl�!2G��n��]Z�����F�QM�C��Ț.���bz"��wLU1�M[W%�`�.�Y�C��	��%$X����|��5�87�\�)�H.�ח����y�uz=1�7�o�ክ�ʉIG9=oS��%[H!y"dW��Cl��,�g��]Ϝ���������՟d� �2ڝ�}*Y'u#�]CXP��e�&���v.����\<W������$�[)@�8m��{�_�oA\�&&=!�꓋��d�ĥ͝��7��o����@�㋜��9C]Hj/<��~~�Fuo�NV���.�x��L��[T!����ׇ�E��o0�OJn,'�7�b�HԸ>\Z�� �?��9kAxV���	q�Pǅ,@X�_�V��h�_��PF��%�}t���:~�>�{��k��ȳs�(�pY��#�2�.'\�J���G��"b��,�A6�'�^�ǂ��wv{ťDs!����l�����	?�r�31�(�� �y�����wm�k!����d��']���?��&q���s@����M�+��k���wD�f����ls=L�F���[ܗ���(���S\����:Zt��Թǹ�˺xzD89E��F Q�fS|���<A�|H�MA��A(J��Rx˄|�΀��2e��]U�ϪS�- ��.ޒ.���8�-
��Ga(�.	��z�L2�Fݸ��<p�av�k�8�O}ľkv����:)2�H����ɣ2���j[1m�U��a�O\ZǄ�}�+��j�%�L]�K��	mY9~��M�q\{�A��o;	�l�`�:�*�ɩ�i�:�rHF|��l����E�;\���R��C�@8e����p��ɼ�p~�K��iW��n�^8}�љ��}^�b��w�����C��T)aM)�Y�kZ��w�"n����A�c���L���/I�;����z������0_M���� �������(	�)��6����ɗ�粪�ViݔőN��~�DW�Sˉg^�c
�x��B�R�bKL�������u�{ы�����W�Ȟ;��R��P�в)K��'hwf�1����t�]�XY����C�^���$ci�zb�G6u�k�.��?�]��U��J�����-D���u������:�����n��O߳�z't���#2�2��+��*V �����0�<�:m��Ґ)�� prRঝl�ܷ���L!����\oV�(U�m�CD��q�#�qXn���Lv�u��D� �yY�2H��6��a/����PTځ�W���X2�U�6�m2.�����^?9&���9X�َ*�@����Er�4$ �(+Ǯ��CV:V|#r�KV�cϭ���}�P��Vd�w_��������)	��V���A�> 
T^k�Q)�	٪�B�{]�.!�53w�͇���%�yzˢ��]S�{���[�>E(�!��2�d�9eԽ�]u0nGz-f�p��t��EZV�c���4)��>�,#UN��0�����F)�Uj2&N��m��tz
cg���x���>� H�W���H;��;T���r�\���p��a�1�}D����=L���.E�@]4� �S	z�7��%�{�E^��b ^�R:�G)(W([���V�P/g9S��*���,#���}$��������ȗu�#.|����QD�<�Lڼ�V��]���I^!��]t��-A�GS�΄k5K��@?��Y3���G��$���=���r|�(�mɕa�C��.^Q�3Noi����Zd�S���>^�8ɢ����;%EF:@�#��t��gO�o7�n`��9���v�:Q���֍q�3=��o�f���>��]��vI���v2I�;<�Q}�<�K�҇�3	���^��r}ه��|���|���i7�1r�y��lC^<z�%��q9�I������'�E��ߏ&>�:��B�7��Oy0ǐ����k����q �K�G�>�N�=�2F�] c�t�
�r����	����Ƕ#v�Pi�9�����=����AS�7S�$Ѩg �c��Y��;�I�f�e�:)6hD�����Ì��T���O[Ę��_��R>�53Y��,L�4�ͨ��c�D%��'�Y����bmN2|隍KA�ϲ��Cy�`��҄�F�S��/��f�nn�<ɑ�$��R��5Pb� p�rg����@�"~��3�ѐ��H8 2�+?��;ji�;v�JD����(7]�pfE�#�K�"��pJ8Ņy
���}��M�$gA��^�$и8{K">�M"�`��C������5*w�;�������XJ�@���a6ۣ�Vb���^�xuH�T���m`���U��8���M�ĎR���M߸�$�0#�xՇ1:\�\��tvŚ	���V&d9�n���c��Y�c���7v-	��#{ez[������<��u#o�<g��tѯ_K:Xu��Y��A�$o��"����h�i#�z	�;̋Ry�$�)�z�����N
�c����)�i1qj "����<��-���)	�1�������M�>o,����#��<�TRG]�I�?!jAS�7E=��!�Lڑgg��au��4�A��W��Â�B<xqa�s{
��k$`h��JZ�7�C;��Fゖ����;�����6�������Q���w���c�3�կs�|���͠�:陑�08ѪڔrWb��F�?2no���Q�{�SxR��=B;R�գ���p�ҏ%b �4 D%���O%�ިg�
�����䏶����I�m,G�|)B�M�_s(J��cJ��HR���F���}d��b�^�H<aw@FR��jQ}8�Y��)2�\ :��
8� �w�l��
e�x[�yD�$��i>���}��mcYDw�2�4�;=��H���X!9�3���
g�o��nN�ĥ� Qq	�5?�>�����u�(ش�ls�?&�Ii�u���`�������[7�G�x�@���B��A�_
�6��KB��x@j&�&�4�B���1C�n�s�+�Mݐ��m��T�P�����-B�x:$��	YXW�3!��g�N��
Ʃ�Q����'��ɧ�:*}Ɂ���AT+�����@���HY��+�+T�1���c�K��v��"}m����ACB��,wl�ҫ�Ըz�k�S�9��<`7V�^l���ZX�:(�,|=t�E$����ďWY:b��Nƚ���8[ѓt
��c����M|�B6�'�JP����~q-M�֢?�hų�t��ﺹ�$�EQ�Zaӿ����$��1��s�h�=�\\w �����v\$��ܪ0�L����lӠ+��.��<DU;f��Bg��M�������D��]��H����y)9�ıܻ���2�J��f�-�'� ��bE�`�>�+���U�&�\� :S/u�rJMu��i������E=ffiwxTr$0��ϴ#N�k��(��������"�2hм�_	f}0B��
�U�Z��9�{?��i|��[�Pe3x�PxA+VQ�C�A�p'Єٶ~Z����EρB�cT�)�r$~���jeG]v�̌g�����%�R��m��0���.6n!5�~#E�����w5�ՇD�t$�*_p�d�3 ;UL��n�����{k�0 n��,g��PSb֜���(T�s3��{��I���Ÿx��W��S��Tǌ���L�`�0WNAЍ�G���$ܻf/-�7�>B;O��=l>&��t���Ϳ�=v{*V\l�+ e�4�$
T%ʂ�,��M�[�b���>���O�u�� �w��'g�%�r�E�DY�ܑ8�Kg��7���]�B�hb(9Aj&��#��;7�6��S[���(����3kłPd�FL�UD����A��������L�QG�ה�¹�͉1�d4���W�J۬nj:���M.�8�n�MHX�|���v����^?C���[�� W��2�^ķ^\���o�~�E�I��᣹�pw��{tY��,&Dq�t�fk�3��'��I�]��kK���h{R���JM�$��N�^[�R�s���#������H�8��'[�,�ڎ�q_:��fٵ�z���z�	�|�^�~T1pa����SPr����Wy}����PǏ@X(T\.�ꬂ�8�`�-�����07��H�|�ÂQ��J�zqQ��Wz� ��d�ҍLqq�@Q/�l�7�io0'��_�ɑ�ۨ�p'�wx�D�❬wB��F�Dc-Y0�F�w�`���N[:�s�Q������f�x#�V�L$��`����f��$̄ �y�D�z���*mŀ9:�8P���oV9j։��W�k����{F��]>=$��,���e�g�֝N�#N�Q}&t.09j-�):�b�!A���^B#߄�D�rƴ]'��9��bc��_2-ެ)�i�(d ����U��6|t�2��60g&���SK��ᇻ=zp�+k6�	�CO��C���8�z��5j9��� ���p���L+��t���`�r�gH���E�q��\ ��-�4���3�i�	�:Qwz��
��57έ��;� ����gR}Qo@��/hK�����.��|1ٰ2��'�o��A�M� ��\�~9b����y��`gg5�X�<@ث���.���X;�zȣ/5���ŷ-}���c\���Il\�I��"��Bq�"��@G�c��QP֘�\]�&4��|G؎	}���;����\��n�������.�]ĭ�,}�KIl.;P�H^�e{�i�(<h_�^mq:������Z��}�K��A���
Q(��v[�& �o� ���C��kЍ��`B�q�����"�J�}#k�($H�����5vg]���qՓ*�esN�iFq�Am�ii�6�`z"���-+a͕���*z<330>[F���K��;N�h~��[��Xe-���Z�""��^�Â�z��2N�s�D!�S��4W��t��Q)R�ر�(F���s����3��
q��b<�ߵ�.�/瘗zw�`1�5w��bm��֔g3�MSg���Y�_�2�ħ����>���=�9Ə�ݨ�E�oid���6�)� ʉ|VX@�<�N!ղ@*zƙH�I�����#�l�X���=�o�硝#z`�`�"�[�(3��б���Q�<���6���Z����������VP���4_lN"t#�@+?Go�!���^�}W����� w_XU�1~���%�,�$�5K���hܐ�[�=C�0�q�q�y��'��&�j0?O��\%S���⵬�4R���]-MG�8��Ţ��q~��h eb�F.q�w��^ı��tW{K3��}Np<l�\F�=wZ�����1�*��F�l��q���	Y&�%��eE%9�OEe�*ּ�[@�B"�6c��"��>l׏�����/�G�ŀQ2cE3�E��BI3?���Ĝ��9��Я������P�e��]c�����8IhʓQ��K�u�̈́&�8rD}?8&�
�-�%X���U���|m���R�u�!#�`���S�9� �Y)(��������x4���QS�BG��f!��>�\�u�	���/�kc�����U'�'O˄�͆bn�x�EPM1���x��&����Z�+��� 2&̓'5K���8�X�mW���T��	Z'��7�4ǃΝ��ӱl�#x�hx���f������h���iT�8�$B_��NI�g�⊎1����(|��2q:oE`��\�ȴr	�J�x�i�Yp�V�z��V�W����g��L�M�#/��;i����,(��J�Ǚ_c����C9����K���] f���t�H;}��Ż��;Ǐ�z.3�Pu�і>Ή��0 u���ޙ��+ack�%UY��%�i5�I�Qj��f@��� _��&�
f$~�6�e� K^Ej�&�'[[�3���1-�8
*���
-�?�'׷�	�Δ��Ԅ�&|�#*6n�P�B��`r�k�R�=
�1�g�� G��1�K��ާ[���B���R�UH���\-�ek�.��M H�W%�J�$��� d�q����D�I�Oa.�h��ю�Y���ʮܐ]ٲ��J#�ʅ�i?�;��:*,��Y�]��w[��V$�{����nvFE�Z��Oжr�
�Ly��
c���Ib��H�M�C�wשi(���O��6��wpq ���w��;��ܜ�{V�#v"ޘ^����=�Y"I��&�i�`���y�i�� K�� �Q?����e���Nb��Z6͆������^7u���ՄJ�`x+����0���:'{6�3����[�Y�Gǜ=�6���I�.���H�?�����^H����@z�����$v��g��U��L4��]!����`�FMj���M���mr��c������)�U��e�� f���
�%'K�-��!q=�1.�N��}W8���O��|�L���8�[.K{�Ji:RsV��Ä�j���N������hju����N�m[��'|-9uV�}PҕO��"v+��)y���li�7l5���'���4�d[�pS|�vj�n
^�5��4����l���е�I�_|�Ń_Q�<"��Xh)�7�@gJ���2p�Gxf� <��*��]8,";1PD��.���w�TĬ�09j��#��$��y�d��)�|ZM�� 8��u}5G�\Q5Q�  �.o����`��Y}���=>Y�+��� !���@
O����E䜁�@"�1	�jj��L�Qt�ÃXrNl'��Hmj\�`����>�;;!I^��Qq��S�m��ko:�Wr�G�K dj�}����#����ޘ<<�u&a�B��3\��F��lp�{|��C�}gC�HH~�^Bl��Sb�Rn�^-&-�,�KyKM�A֕��R|��]w����㸇6�J0�T�U�I���1��������2Ȕ3蹧���~=Rv��Գ%��վ�Y^Y�Jk<��4�	��-2�[HDV�$Xk�#�qdwڈf{@�el"߁-�(�/L���Մdsم!òf�س��@�����P�9��VGV�h�ux��M������\��VU�,Y�]�ssM�FK�Tg)d͢��L֮>��N���Ӓts�*����a�!� b8��Y&��,2`,�|��V�A��ѱR�8���T��̹���+PA	9��g𳐦rn�n���ίU�V��ll���������%�/�x���x:��������}��i��1-� ���q��st&�gZk���~��E��>�CP���Ne���5v��Dw7oh��̼�8�}/b���%�R�<W,7�a/���1O����^�7R�h/�ΨN�5�����(i�}L3�n�)!9�,��֣R����z@��ݦ�#E/G<*�+�0:����^$s��.%h���Ug�:u�S=U+�F��9g�Bn�ljHa�斀ͺ@XqS���I�c��U��8�1����G���yu�V<�W�"w�0�	Dh��8N5������+� J&�R��:?<woN��e7g�@�f�Ǝ��G)Ӏ�T�DkRi�~��m�s��I��"W�b���<�
��vs���ڥ� t��
�/qB��r�q�73�O��������u�g� ��Go� }����D��#�*���c ��A��\�`<��c��N���ʙ��
6_K�'�<%B�#�\	7���붮�D��A}�ݖg��Z0ϬkR�F��/ί�oYA���w�0�0G�)�oh��m!cW�_�Zq/���IxPHhof0����򰪏������O���;�SKt��A�I�^*&u��G�S۔�`���x�b�E�Q\���H�,Q��+�m�1[��*��P����#��>D	�\:ӕ:l�O��v%��f���0g0e�he<�D���	~h�U�o��t%m>7��l���N7c��&��8��"(�]�ǐ���pܷ?�~������?�K4�����[�ۤ�j�6�&4G޶[����l��`��`�q'���!� �6�vi��p�����,�i��z	����AQJH� H̸�cJV�˱'H|rA��_�tp�po`�DK�c�STpc�
���A�{E�:#�!�G��N�f�=�v댞oܒuxX�����_��xH%w�� ���E=p�Ϭ8�:�\f$tM���e~�c�{�g%)�E�b�8�%8Z�s�K2�i�'g�VOW 6v�{5"�%������~���a�ڙJ4�ri[��?1�`,�ŵ�y,Ĉi��ET~5d���n�~�x^n� /���^��ɤ�`��y����h��S٩��Q}�F�.{�ԫi�|R��>J��{:J�m��]�>ܡ�4��Yr��[����/�9��6���|��?{��1�WlI��\4H��4d��oW	J��*����B�($�V_�dF�l;���Ot���սu���T��~�� �:b���Ʒ�����*`�ϗ�\�W���d�[Q��� �*�ũ{�������`�A���02O���M�U�N1�ߚ�֞�ה���� �+]�3�]*���t���8V�o�͒,�t���� v�"�BFYT���ڭ��Gń_I�p��)��0���I�RȽW� 1�s�����@�$T�9Ӧ����e�@�&��"��P,��e����Q��$o��r�����I4҇:�E���gέ�+I1m{p ��|�Թ�LGo�����@���L�+�Wuu�J[���0e�m]/��O�ehv�\GPB���=č^��b���q�Z/����k[���uX.�1���<�7v#�cc�q�ɵ�'z������^Bzm^��DX�s�������)���:�E�i�H2)k���t����ijC�X�r,�Vk4'�ʛ�Q�5������0���x���K�ACp�ى��oo���q�-F+"@ڡx�![�c(e�D����c����$9^�W�i��������l܍ѱ��s���4�1�`A���ƶ�
xL������1V[EUG�����>$#�_-I��1�31�����a�K��A^�-��':` Z�&<��f���wC���Ӷ*����|�ŏF\B���s�D����$$�n"s�>A[�l>k�9 a��ӆ'�t�+�F`XJ�|QK�xq,EI���/T�bq�@&�k1��x�NuԎ�h���97��E�]�'CI#���,��mN��=���M��>��|k?�:J?����OB�-��Uo3�ԛQ�/cS�V����rÀUgO��~����#�R�ؔ�8L�⣥���8[����?�:��0�Ws��)/-��Bч���%��eHH@�Å\t!�%~�#s�,f�����4��M�ò`���{��nm��)-SM;5	�o��j�H���4Z�mjy�1���,x�"�n��^/��v68&�������!u��L����Xnj��8�+�+�ｓ��o�����JX�Z����Fdݺ�(zޯ}�q�&C�-na&e�.�I[A�!���?/�<�O��/䨒?@r�&<S���
x��]��Rd�
ݵ��n��-���h�^�ܙͲ[��b���;wZ���=s,�=�f���CݍbM��|�Tӆ��@z�/7 �� �۳2\9r'�$�b:hrr�X���x3�(�'.I��������4��y�fgU��8��2/�{�K7i�Wʺa�n����y���$5&.� �Q��������vj��R>Wf'ٍOR�~&�.)f �-�x
��Gc�&�|��#h�w#��_q�$��2�.�ۙ׵���O? <ڵ�T�u����_m�O����}�b�0g��$�<�?�Ϊ�>�,G�|�G^��K4��$�1��p}�=7��X�Q�߂���W�TnE$��k�E���
dd�Ek!r�X�����@�,��rė�[���M�(�� �4�y���Fj=��O��rB�d�n��
��\�c�8�H:��ja �GH8�f��0����њΈ:�~[_D��	Rqu����,AX��x�Msۨ��o�R}`˭�e!���gwdW,�i\��r��=�ua�	��c��������-�X���NzzT�j�Ae�dֶ%v3m��5-���0[nׁ�_���B��Ad#�k
Ӯ^��>/��g,�'�	��2�K��
xP����n��̦����(��o�;8H3��s �knԮK�u�tIC;���op�v� ��z��P����u,l�tt$8�=/�+��)���X�>31N8Qo:�o^��������2�h��Z��WW�����[�a�;�S�8�Ǯ�"cʎ���R�z*��mKp���%�%��WѶC����sr)�E���=\���y�`����ʨ��O��=��z�(jH�'�KElK�0�hm3"�}%���)_�����6��N�Ӫky�tX����Q�>�p_gqWy��
#��D�ں9�{=�,(��ibf��5�b��a��x	f
�������gʾ�����[�w�F���Ӹ��w!5Q�5�t�B�X����d�]ٙ�%8����ҒZM I-Ӡݴ=y�9��jR�R�E�� ����8���do8PCw�H���;�,�ŀ���}-d�z�<�B>Y!����g@��q�o��މ�ȷ �n�2�� wwW��t�
�T��"k0�?�#rI?|o�=�,�}��B0|74A�R��
'�ޣ�z�W1M\��g3�x&Kb.�F!��[�A̦FH�����H�����&¦ZF�7��A�=l�n�<�Ek����r+:���hH�81nKv���Ts�j}u�T]2o/%�=
�E�{3�0�ӌD`+������5X�j�4BMO��1wIiC�Q�~=2��q��j�:=�OE�o���I����%��;�3��$�3��N�P��?_�{s�^�)�)���m�he�8��D��	��^����U����`�]��ߐ?V�x��#s'��Es���b?�Y`FK'����_�!+Oh��mFsMim�����y����V8:G��-����$4�1���"U���	kl
�"�)2)�����#4�7�K�6Y�U�m��`�ǻl@_CC��`�m���<2z��D�+|��y�����D�_=P��´��/w�:(���
�����j�ٮ��u1��S�����M��s� �茪\ l#N@(�7	��xH��&텡�)_U\��N��}�9��[� ),�F�M�9hX_k;w�n�~����G�T~\��d�,`5��"\�L��1_v�T%���_��P`��_���<��O������a}��&^�*�Ӈ�?�;IXʃ��;�����l�������#f�=�wE��9���y�_%�#�}MF�h�{^F�R0��d�S��lS�@E�2��%X�3��pLX`�h��%U�m���t��*\�CO<�@T�~�̏�$�h���Q�'+RH�]G �9T�>��5�m8�u��-���4�TB3��%�s�3R�y�2��B]�ՆӍ߂-����&��}ɪ;��!b&�R�}-�i�n$]����΁!���D5׾�J��<��z��c�{t��sq����׹8^��g�u0J��\�B|Y'PЧh�z�N]��� J��C�es����q�n_`.y�l;������U�!���yH4��Ʉ��Q��������R�Y�<�. ϫ�_��o�Y���|�!�`����,�.l�v���7(^@a��c�ہU7g��-a
��)h-vy�d6-u]�u�
϶.X�nrҒ������h�5+�:����#�պ�&�L���
>���V�����	B��c�Ƴ>�/L��-	;��A�
Ԣ)GD��L��&c�S�Ʌ�l�̙�å��x!2�PAkvs�s[Hρ�5l/%�:���XH����Qi_�6�\΃�ɠ�HIX(�m���XS�6HU���pã�ej�	�)t�u�J�9��7���`��g��D��-��+�=��k��� \q�E�(��!����I8 T��@���GlO��v�&�W��_��A@�N^��D�uqW�Mg=����2m��*Y-�J�9���eF%*����Ĥ�@Ϝ<�y�N?xqi�t;mt.����E��7�Ar/2�Vy�����/� f�0�C�}�Wh�f�F�b�F'ɯ�ռ~���t�6�������ߐ��G�lw�Gu����*�����x���� �\Jv[y���4���Z�/����Lg@}>�lb\J� �"��/w�V�4D�+Z� `N�{���Ұn��{^�I�0�2� ��&|o�w6\�gX��"������ۚ�4�ڰ�I�Qn
bq���!%N䑓"��Mk@l%� �Nm�����x��N:�
@��ͫ�e�*��ń�6�M�2Io�Vr�
'J���J���r��pH�c��oy\�=0�������_2eW0�T̩���$��Y���5��+�o�1Q.9���[�.W�Dp)�d�/.���(:+۾�F����uY�T�
��
��{ʒ����*�[�3�)��t�>~�-g���N��nϡ]�,'P����,E�y��4C`�lH����i����cG�p�ŐH+.NU�D:����Z� e������o�2�]Đ��1��?�(���^?ys��[C���>$���ĉ��$uT���7fA��$�6e����S�&�p��E��L�$��	Td	�7#��r��hL�t�Ƞt`�xF٭��F�Á�]tk�Vz����V\צ|��\��{Z��Z3��S��L\��3�X��>?F��WS����å����{<|8�h��m���0����ӽ|�J��0+�-�`�'2xXc���"Wr��k��T�H"ŹF�ǅr`�sʢ�:��EŢ����^w.�=�a\~~J�[���8��/4ɀ�$y0�T���
����ȧfD<)8��#�o���W���k�s��!��_oz��M.��ʂ�wzZR��]lD���@�^L��w�,�a�6�ӏ��F���/�Վ�����2oZ��
q�~,�a.zE���
ͮ�r,@�sx�gk��a!���3/��9u"I�w��\> ��L:�t���D<��\zX�'*<�SS�w�lҐ��8l�~�߾j7f �Ra<oi�g���U����g�|��pGhKw)��(�4�#�GYS4ّ>쾩.nJ)�e*��!�>R4��J����p?C��kꜴ�Z-R���x��h��#���M�B?9]�)`6!�[7���w՜g�ym�!	�r��u�x�B�>��^�;Y}����,��R�jV7n��Q�2������5?+a�a�c �zP*�����tJ���0s޴]�>X���Vqc����e�cM��������� .F������������Wk�6�W���o���\��3�$��4���U���z��O��M<�ۜ�
��ɸ�?�A�`(�&2�K�2�LF�ND�x�n��T�A�O���NL�G�3n����#�_��uNn�<�\A}^�kv�$	��^���dP9b�7uՃ��Ep���f짐�K����K#qem[W0��F�	r���]�B��Z�T�=��[�y����NO%U���D���,&�����Cz	�cx�夽��<V�TSf�����o〲�l,.p�� t���T��hn}�*���'	�7��L��k��xM{���k��Ӎ"0�`;���g�Lb9g�'?�5��nX\b�Pj0�́�~^ۨCd�U�.؎�a�F�/>���$��!c�����8��g�1
Д�p���x��� Jп3�K��a.@�՝U�5
��E��ġ?SZX�A(�u�g�Ë���I[�M �`C�& �%�;�%�\����;9�I�yyt�h��#��<|����l�L|��~>^.���m'�us 4`�p( z4��&L���\$�%Y����ULK�.�3��'֏�( U�IM`��j"�f�y�c���d�#�u�y�w���������+����|[|�?����GЛO%��W�OM�u��1l��釣�:d�%��yF�,*��(em5�%��1j.mp#���b�i7ն>Z�6U&�.L��.$0�씐��
��k$`=�ɼϠE tʻ��à��ķK��a
��*��Ee�����i�Er����y����O�#���4&F~��v���"��k*ۖRt�������`���Hm�^s���A��%���\2
,V k�H��l��� ?6�zfUO4��h����OWo��wn��;�o��/�C��e�������d�y��4��|B��xG��p� �rg ����� |�<����*��A���,�>�{^N��͒�Jz�0���%�O5�x/A`=�c7��YZL�W�:�J����(��Ń,8g{�aKm>���l��ʏ7}�E��q�4��O�mB�����tA�q<�u���[2ק��a���� ������#�o@��<T؝���P5��6JC�ɫ��Y:�U�˙m�˃�uO/�Z�q�[`Yۈ������N���Gg��Q����̊/+ʭ	����w��ծ�MiՖ\C���^�R <�I�1�����w;�4qB����VTF����~f?�q��~5��B���ފgž{^�����,��ۦh������7()y�-z�.m1��!��~p�N�g���H��e�i�0����5��X�a�=	��3ц��Kì�����3�Λ���x|�^/w��htH$x�Ō�F@6�z�_أ�?���,���ԁIQ��z�h(��O'b�L��L��t��:4�
Ղb8��2|�v��}|�c{a����W���w�1w2�L���L��헟ou��:F�8I���n�+�%��uU��]C��~�����ƿ�J�z�o��Х
u��py \�p����v�ˁ~���a|oA�;�mrԆ_��E58�0	ې�oDv�Q\X��nG֞�|C�����z�dPT'Bd�D�2W ��8��lPD�Q�V�$ITω���JM|5 ��Y�E��%7oԖ> :�6��#Չ<s6Z����m&[-��b��ѝ�S���נ�gC��f��������V���xz���b�%۩�`�̺�;�f���Α$�l	k��ȇ�A�ۄt'6w0n�� �S�E��W}�پW�1HD�!U��Yn�
��hm����-ؔ]�`D*�)�9�]c~4�w���K��O��r�:���G�4���l��'w����/9�JPy��aza )�J�z������~X/��D#��_E�b��;���^�����o$r���Ŗ� b����b���bb5Jl�[��Ї���k�i�*�i�=�;��7� M1*S��R�)d����˱���D�.at*������^/�{1\PL�]��
.i��$��`"mx������i�Af*�]�U�����{k����qg����Ⱦ)#Y�D�߁�ml�^θ��dX�]8򣋹�RT�&KV��^1��&��e�̊1O�gH�Pn��[�K�i�����M�B.>�4�`�L�ګ�l�9�������S���f$s�w�=���Ԕd�F~�8_$��f��l�2�*��`�h���f�/|�I$m���{j!�8<N5j���%R��bAc����$֙���x�����*��f�S�	��B���ٌY�sk�Z����3�'u��E����vRL]-s���o�y���@}� e��E��gܟ��h����A'h.��`_��Y3U���b�0 ��Tի����f�0LEU�����<���T���W�Y����*�K�U�-2�39sC������K��V��c{�d8������a �Q.Ѫ�J��f; �4�Ы�6<��3�/�@T�/��l�
�Z0fγ�����z�3����H3�Wbe�Z�!ú��*E��2��֒�0�b�M<<6f�Ma��*���*]��瑱��:�)�Jj�<eslX8��h��!!u@F'qa�#g�֔��L01�A�޻ׁۙ�#@.Ј��#�h a�Ԡ���y$FQ�t��\8V@MX�,��=?��$��,�Kx��R�r�Gb[�򸮚 ���$k�q���gB� ����`�9��ܻ�'/0���$�|��35oۺ��^����Č���a\u� �*)�u܂��K��և����ŧHȧ#�uӽ��lv�^/.�b?v�*#Y��䧑x��Y):v�)U���\����.ж�oY���� ̃d�VAq��D|X������g�h1��wWC��Pߴ'e$ SI}E.�#�|��Z�ʨ��� �M��a���.ʩy�,�4|��u��?���E�������U��k�J,�z,Hh
_�FPI����L'ީ���e>�����?N@4Ʈ�4���Kq�(69*ȵ3���xH��]�@�ɪp��՟E��js!�u.V�͹�`	LB���:>Zi)�y_���k�/����җ	#���4@���Ҷk�,�H����xg��������L�v)�f��M���1�n���C|l"�3N��:�j�P�=���d��q���ZDf2��N�av:�n� 	Z�_=�X|�O9���ѷ����כqw��m�3؝��z!��#�����0,�p,,�z�
��b ��Ġ�6����B�t�M�����0"�ꓢ0��`Ե��~��><����G���E&��l����i�����òF����+�Yʺ)����\5�>^�	  t��z�A�e{�J}Ʌ���&=j���.�X������>��h�08+��z�A�u5F3�=��Q�C'D;���[���8"b��F�׸�P��K��-P� ���zl"z�UA��3wK�lٽk@�V���hԴ���a	��_��a l\��pvі|�,5�#�c��tYJl�zҾ#0[n�M��ͻ��ҸJ���i���;��v�u
:D�Y��i���Y�rp�6�Y �j��A[�P/z����Uu���S���7�@�b��/9��o����I'��Ks%L���
K;,��BA�W�_W�R$�g_J��q�f[x�m���7=�g�GZ	_��	���t��b2~3D�l#�UL�⸗��d¸�$�<�;�Q>�l���u4��Z_�-����?܇�%�ȍ7\��__,��&�ҵ�Ǽ _|�_`�o�bR���]^t���M$/9
�����ۋv���"DG{4Z�#x��S��_ar��Z��4� ��\��. �����F䖰rZݯ ��By�D�6xO6�&r_N[�e,�q��j!���4�V4bAza��Z	BV�L�7/�&7�z�ڹ���\�O�%���3��ޭ��u�O��	���N_�����.�!i�G���đx��QujJW�����D��U�ͩpl|��[�H/M�%��{�of���>P��ȉ������x�s�#�$��l���x)X��d����Z�s��Û��i�y��$���<�O��Lpg1	D;�R?\�hp�B��T�x��M��u�8����#��(E<u�ͽ�=Au���\-��0Q����k!^�������J�G��M�g���3@�h�O�d6Y@�
 <$?f��|�������F�mpnt +���-_ЧF/g��)�b'o��X\f���R �ab1_uLJr��y��H9�E���	zQ�~QD��w�S]�v@�~��b#�l#m�Чi�{�4*���.�M]�x��}��	F[���~T Y�;���j�+��k�.��3¡8$f1���S��f2ՠa���/�3P�	G#����U�[��t��4'��\7���mXh�~�E�#`�>�A����!^z�� �s����1`+ԭ��;�/V��C��ĝ��%�Xo�ng��m������]��n�(�t�k��&�,�8!ĿjͲ�D�}U!!_cv��PYB&e�V3�䒇������Vd�̤]�e�ˀ���g�@"S`�# cս=�
�,P@й-�ms�A��5p��2�&��!�`����D���*��}<P��g(�P'eU5Y�2���*��}{��.����Ǔ��,�e�U7������籙EO"eu�4	�dQ��3:��x����Q��YE�U�[�"�e�B���t�l�1]�*T�bDi�S��CMx���jI�PQ'��02�4 6GF�Y��V,X.5Ǝ��ć��qG�A�����c�ֆc'h�����R��]�������v�^d��?���4�����^ ⟫��weNd4��;Ē�c��{ql`}N�ϘR�Y�il�ʡ?LY�gKAZ�]_�9?D��K���k��Hvt-�]㨒qy���'�;�G�.���]g���������+�Ҩv�:z(A+7p��{p�MƤ)���9��S��uǺ��R�  ����A7�e��u���ye���aF�dZ��p�!z�$�e��ךE�`�8@�l��z��mf��mHʏ�Ow�y�tJ*�4W�uN:�t��5�dd@۹i.
*�Ǳ`T��7�,��-�z��d�h�HG��%=���'�5޽�\|���o�ވ��fuk�
�E�R��Kl��I=� �ʔ %���$��wŋ����h=��\Yl���	3G��B����^Tu��5.���$�׿'=j���?;��h��V�\5�������tR�ia��N<��L���xK�Y�B*���[e8��!��*P^�%O�����������i�2���Q�Vm$Ebq"�$�p�B�U/W��zN�/�����,�q�^/���i�@���d�^��u�󇊭�����>���]�C��(�H� Ƒ�01?g؅�aU���#X�:h�i�D�k�G$��t���nT�#IɁtN�6�3:���F�B@嫝���)P)�e�埳׻]	jF��cd�$���η�J�ڳ��Fk�{��cķY�.�w_g-��]{g��|��i,�PO������@~`�f�^�B:jP��cT��Nl3O���OY�=6�~_q҃w�JV|:� R��v��p2e�P��Q�a����>��o��H����/.��ռ����-�}U�s: �O���?QbB=�g�1�%�&�hA�,�20��by�d�ܻ �|����=����;Y��Ut ���O��]x�k���ᾃa�YE�:�b��h\-���To�B�{ϵ�bl�[�A`��5���I��hZ��>HW�}�
���EL���F��g��~���`��>�2�W��b`��N���Z�����b*��uOc��
d�$s��
����(�G��OW��H�!*c�̟L@��q�Vl������A��1�X8Z8��(/@��ff��3w�K:�<5\�t�⪲��g%	�S78��z�޷pt�G�g���*�HyB�q�,gzU����@��?�h�)���(�]ԉĩҗTF���c�k�L�����>�:����'�Z����Y�3�|v�P�F��aF�#���V�z�ją��Zt���Z���F�Y��`a��[�|�緰��i������,�ham�b&7���b'&���fRI���7%^���Ԥ؍k4�Rb���[g�̎O�Z�O��k�����-�13\�Ǩ����1�7�b>M����/&��>��8)X�V�q:�J�??��P���+��0@d�}�i��1�}�.��
@���	��9��6j���pʧہ�}Cޮ2�wh��!lc���(�M?A�?r��9�+��'���n@�y��.Ce�B,6u[gܽK4g��WCloA�jzh�7i�E�u��_C���Po�<��s��y(�vj���p1՚$�R{�P鶅��'a�_���@����f.��փ !Ϭ�h����7E��I���m��2�87��"jcF�	�[;��	i2n4�C�b���%��q��#w�#�
�[D�k|��P���%��VS�DX�u��o{}*�� 3�Br�
1�`F�g)M���`ֳ�J=	�"�ND�����1o���|���T��!~�'D���r&LhVLn1V%��{���1H�wj�8'&�8��aB ��{����[��Z���a�5��0Z������o-�����%ԖU_�
�.�G��%��X]S�D?�`&�7�/ �^�o۵�-mq��_ +,Cٳ�#�F�N��\\$�,{�5��D�&�;	�{�Uk�#�����?���ʅ6O�+C�4��I���1� ��α,Tc��ȭ�A��23L��y79�[%Oe�>�q��r�X/GV�/�����D�.M E�k��4�_��t�F֊��G��m�(^8:Z��fs�0G��Ă�I<0Y
ݒ(�����a�(��{��'��^�>�&�EI��1|}���m�����9J��äę�9K���&��V~k�WԷ�>Xo���Yܻ�G�����Q5�Ӛ�`��P� ��Wl;�)���5��-�.��B�ԯ�o�(�Zq/����(S]EǛ(���SvSLX��h��G�R��nP�7��$K�֪w�u���m�[���`?-)��3@�\G�n�b���욤�k�5j��o��-�;��)N��8���M��J�4������X[������mu�N���.���t��~m�n�2i�b3�a,��ٰ���8T$���ٰ����3w���f�-b߿��:�e܁��c��KȰ���C��@����蝒I�L?� �E4��/'?���O�y��0%N
������qxu�Z�^��*�K&�ܣ��u��$^ĉ��Eɹn���?ar�O!�CKe,��U����ḳ���X�8�\�y\~����c�u~"i<ˋ�%Y�X4�>��@��|�ǪB\���)C/��K��2�*�8�:/qҼ'��.|^�w2׀x`�r}��4���.�@x��6�/�����&^8�f$�n�7x!ԟ�K$Qy�k��C)[׹y=�O'���P0�'^A�p+TV��]��/zTb0U�si#�'ec��d��PѬ�u�"k��}ɗq*uu��M�:; '��^dt�����ɏ� �,#�Ӌ�T`bB����HĶӓ�X���3֫������K�V��6)6ݐnl��:����D���e�%��M�L䷜�R�%�s$�N
�r�������~�������[ptC���
�f_o���$��q�'����8���2�G�f�q��l�d�N|w��ِD�9�������]ڕϨ|(�_U�ѣ�+/�}��=�~��l%zF|ѹ�K?�0��4��H��j�4{$&����E�^~SR_D	^��*hz�ki������i5!|�j
4`@��p,f�>�A�r��xݷۤ��6N�a���z���iq��H�p�$M�-��r]��3^*��>vD ���s�fL',�V%K�q�Y"�Z����= ]����&0k�h
�8n0��W��
��w,[v�M�n~-��*JA��b�o�^�2J>���*%�+��P3��ؗ�v���1���~���>ը����0O����6��ug[cI�=���>]��6�6ݭD�n���E�p>�ʅ-7��t�A�������zLǱ�]	�X�c&\j���h�1�-Y5D��6�R1�D"����) V�g�6��Y�D6�#���hν�Җ\%��s��l#y|��O��2w'�fHض�|y��0J[ǲf�[�H�JK���E�D3���*A����	�K�(�ց#����P��!IٌܫՕ<rWl��*�>���~.�����@�I��1��êS.I
{���[Y���5��۫�Ҁ���m�� ���,|�_�)�G`6�Tj�������.-���G��M��������s��gr_[�ԳR��h��P�e�Y����*��a@[ޝ��%Ã�ӄ��#>�d��;� :e�16+g(��ӴS)�|�wB:)�Hǎ��H�����[i�lzܬ\���6U
�Z��P,�L�?��e�+�2��� �&����:���L�����Ǵ�8f����>~�1���-�����È��Q$����v��L8���=��@ <,�!C�O���|iӽY(��Ŷ*Hw�ٜ�>{N�q?�=\]�4P������4��+���/�1��n8��,4�8�&I����ڀ{���s@�[�@8��T�y���k��C�m��ix4����R�,�Y:��}�R��y��&�=��;xK�/�K�T�ɫ�r��۾ީ�\���S[��GY���*yhd�=�'@�g�-� 8�C��V���ժ�3��)��z߲��c:*��-�5r�
8�@��W��-J�ퟥt!�g�\�"�2"*����?��2�-���-3���|Ƌj�
�0���d#�(� Gȳ�F��b�Ho#x>Zm���Ah���B{�H?�v�a�t_�+Ҧ$w�\	��72O����-�	TW�[G�������9��H��eX�Њɼ�d\�
��sPMxY���J�S�붆~��zv�b�̬���ڹV�~d:m|Jo�6���$���	�?g�q������WB�rc#H'�5�P$ԑ9t����t�h8�G�ߛR�=Q
0���&�-�%�ؗ���a�$�������x��:�	�+������Z
��c`#���%h��AdV<9O��w�e�<$a8�P�Y�u�3��Ww���V��9�wr��3*Vi~Ε�d 9��`���/�:BE�۞ɵK��0Ƽ�,IU�JWhm�_j/"[Q��ޭm�ͧh��=�u��a�O�蔺�&�X�k�D��#B�r���%�~���%�����2CJ�+��n��]75�pC���KM$�Vo��z���N��v�2&��϶տ$��;
����v�u2�g_P��M)���s���Z�V
΍3�;�i��"'�S����Dj�C��_a:A���^���q�	z�~�f�j/"r+7F,-+�R��"7�Pr���r�`Ͼ���s���z#W����Q���c����%̫~߿�x��!��(���V�*P�S���i�@_"�|>*��JřHN
����d::7|R��h⒕8zY�M�HH(Jgה�ޝ-��.$M��eh��B�SRՐ��Lx�ۢν�x�9跕9ε�����\-Bه���v/S�����Ԙ�'c������1��ި�I�$'�ۻ��.���<�-�{����;A	�+-څ�1�lQ{���r��U��2�߼,]ϙ���s�1D�L���|`�.��w�`WB�#�#��Ū?37����D�w�%�v�ye*y0�Gz%����@�b˸��/�bx�~}r[n�L�E{��V��l�ĺv�1��9'���	�S�5�3*�ta�q�f̾ �8"��.�к&D�w*o�y���]��k�=>i�=��G����O������4b"{p4&��p,S������gA�U,>�:�3���%�9w�тE���'�cp�Z�����a��Ѐş
A`�Z��4 
��wg�{��*̐��r���=������yƢ�8��uͣ�?z�ORhC�V\֓I�P}c~#��Qd`ήfD?o��_��Y�^0��5�v�[-א�wU�
h�ٻ����lo7���Z�9�WA�Њ޻�g�y�<5->$����ݧ���V���v^��	�7Ň���w��q�r5D�da ��.�ݼZ���f��AL���]��m�{QL�U����`�^��x/h��c
�ps�Q��;��6�g�.���X�+'L�}G㗂f�}�#�M �w�x��I�̼��G�.E��&-�)�B�q����!��l����XuD�9aք�
8`��:v��e�! v�έ��q�Z��R\���G��q�چH�*�H�
�RF�[�\"��Mń�%%�Ё(imp��YG�j&H�5�nrD�B�A��u�>+]ug^pQ��3/�2�Yx˜Х�����^ê�v�^�w�_w��t�}��и��.�q��,_q)cA�ח#��eS��z�{xӏG���QUڑQ�؝�q�3Z}�9Y�A�`$$�d.g����Y6G��J�YsCF(" t֛y����=�J�b1�lԏ�T�d~����009*�/���߱��ۈ���c���󛏞t�IQ�F�Vɔ���|�Ox"���@�p��0�$R�.�7��~c����+5 ��@�ҡx����\��or��B���`�"��/Q��ԅ�cZչ��rG*Ά�\-�~V9�Ų��/���FD��Q�� ��0R��҃w�8���$x�Jr���J��t�o���9��_>��Ĺm�0�9�L&(��1�Uy�*�K�ԎK�� 4zz	�5Z����*r,G��6t�69��8�����r�&3&���j� ��K���a��@�eJ�S�䞋����Wc�3�+�%���S�_�<�Ǔ�y��#�PNxx�{�ie{��ax%U��ۿl^�����]�w���b�|o˄%󒆘KW1�,����y���JYQ��:9��j��Ӵ��>�M�B̕)�6&}�#���Q��ev|PZH�wE�U@�/�!3���)�� ��.���y�!���Q�QZ��I�[|醊.��2^��5��ua]�ί����n��f�]g�����vaE+���Pˎ�;���f�Eחe8l!/��<��=��y���Py$�T�CN�� ��� ����qbK����d��C{�6�f�-[-&�?����Av{�ϩ˶rm��~�����)>������a7&$� �̧"�&�����.M�-�ZX��-�c��S��o0ip��0�B��G�g�&�[�!5��� ѫK�"�e�u}q�q@���<2��g�O?yz��v]���8�6V����q�
ǄH�u%Ȭ������'�]Iv^�@)�/z�E�w��n
27�5َ�&f�N̺!N���c���7w�Lh�4P�'�D�Ąn6�#�`->yMw>���D}����g�.Pen���/�Z�T��_�n������;
%z�Fj�3e��e�.��V�F6O?�7�6��.':�A��L�$����AԞp-��]���K�o���'Ǯ�*��뮼C,��K�����d��r<�ߪey��!�uW2g���"�$�F��*�d��D�M�-s|��M�W�Oh[�ҮH
V�g�B�j�=�4���y.y�feC���fX�g�n�F�>�h�`t_9�|{zk2�ǳ���a���W�ٮ��5waX�L����f�1�%�����zDY뮞4C�*CC�9Ed�%�l����,˾v
�\s����lR��T�w]���0$S`ߚ]oq�nU7ظ�pQ ��M2z>�_�"i��XFg�[�OM�i��X���1��6��Ǵރ�>2k�4qh���mw�A��〼f.
c
+c"�ʬi��r�0b��s����I '��|�1�;`p�ʍ�?������E=�A�� >�F��Nw�I�]n8J@
)�)zYw��߱Jx��ϒ��e�ڢ�'L�v3Y��k<}ȷ�=�7�Ѡ�~����	s���>�;[,�7/��`l��H�h%؆!m��}u�D�I�(G=�ST
=��=鏥E^*]��we���������8��ʘ���Β��`Y����/F��(��XH���3E�l��<����fE���:��	Ǉ*֭e8���D(�𨃆-t�x�[�_��ڻX��� X�ɚ�=Oƽ堿�X����5��8y��i<���A �j�-z\�������J���V�vu����T�"�F�t������T]��~�WO�Z�OdW�on&c�d.��q�W�"�s?#ϓ�U$�q�o�� �_�
aԵ��,^z��ިj$��Ӝ���I�F���Z,�&��E��p	|b!�nz\G�x���z��A�B0����}�Po���
�V�T�T9=�S�qV�-��9�.I�rȎ>ꉴ`
9����X�=����U��Q�và�/Yحkh��aW����w�ï�vI��ۇ�p�G��ة��J,�	]k�)�(���,��/�����W���Z�w��#�g#�L�!�K�ҞU�A[�7.�ǐH�`K�FZ^U��J���h�U8J:Č������!-�jB����K�4��
	Ur/4���5��k)!�d�JV����>E�->ρ�I4�j�P�M���ؾޕ)=�`����5�{=�q%xx�ީ�aq;K�(X7"��c�?�%��lH�>^TL>��5�H�]S^�W��mt�$��@mF�>ahI�ѵ��E4��+z�@�D����J�L�,��ar��N�r�n�����=�[��q�����֊d`����j6�?/
g�jAI�
�5`�G��6�P�D0��F�޴�-����Wn�{�*�ӻ7`��o�"�w�?��p
�)O05ns.�Y��CS9ǁO� ��D� ���@�އ}��/Ҁ����*m���-��U��V����:�UMh�n�b@�t�;B!����y�"u�%��e_%�u()�&��l����Su�qv<[������8%Ek�d��Y���嗽6v�jy3��.��� �j�vQ0�e���̋��Z��D������UEI�F����=K��D�G��(�@�?����|�?�Ϲ;TbT���mB<!-}nN�=딣��\��g��a�����f`����%���=?Ƃ��gV��Bl}�a}�~��\W����<�j��;��qBM��^�6�>�ԇ��v�僦�i�|�����0��S��;�Ou���*�������ʬ����]�y�tN���9�LD�[�6������v�yu���5!�k�t�g�;��6,�22���ߓ��,,�{q�������N���Q'z�n�Ⱦ���
��.����㐉/���%�d��U�׳���~Ꜭ7s(t�E��'`�|�A�`�8Բŕ�\'�q�v��g�OBʄ>��ƿ�5�m�Ń܎�[dfi��	�r���{BW����%~s�C���I����W�n�|����B-t�l�U��(�����o�>�a�#���2}�:E\���0n�/y��\=��UY��"'�U�]+��s�ݶ8��p,���%�h�X`�H4�+tP�B=K��c�%X {PԸ���TO�ֆ:�^G'�f��2Z�? �p*�j���KZ�,0'<�\�:�m	�p��w~�.z�nF9+�#�M�,�\�x� �*�G�f��w�TP2�Z�	�#���n����$;3ǯ�W�j�5L#٨�/�h*/�
r�4UT�������=Ă�po{؃gجs�� Mv�����R�3? ����z���,���U}�;�,n= �c�_�0׉���P���޽�P�U�peݣǋ�O�+��=a��ї����f��T�����n��I��Z8q�T���3��
�$��h�(4�%A��_z�@�;�p�raP|�nu�]2}Sp�x��&���tq�F/3�S9���+D��E��Zt+Z)��)�=��׶��&Yo�]�������:7������űv͏���g�(��� �P�W�����`��ㅅ�0�
�]�[�Y2Hs,�� �M�������p�/
��d��$�A v/a@�^�ab����;�\���&:\'�t��`��t�_�=���j�p{�P��<l< |�k"c���s�lZ�]�Dr��V�Z�&z#�Tx<���� �~4a=�YF'���<8gY}���#L��Ytq
�	R/�O���,��*#�}i*���\�������5i���ʽ�=�?�x�����k��˶�λ�~f���Z��&���m�7qN��
d�d�ر���{,�ݒ�h��H����f���kll[^�"v�Y��yH�e�]�1�&Ҩ?X�)���ҟ��#�� ;J��mvn���y3�8݃��R(~�(��
-��8��*j,&C��g�'��� �%Y������ ��������p�n��-k�E2�_0��$��#ɝJ���q�����c�(`^�n���F=1�̨aa?��$�w2�="E�X�$����,�A;���y��K���mC �p�VuZ%�V]2��!̣Ğ�d|q��i�J|��Q��׵'�{��!5���� �J�^��Җ�����3�;��S��0�4Vc���9���&�w����#���+!�!t��Sf��1���³N{Ik�Ƈ�.ْ!�.^U��������Kf�%��tn5���%ЦĤbj�-�����ݖ�\�tf�,ϣJ��7p��I�W3ԡщT����R�<�u���̼ZwL�l	��)<y����g�lܘ`��� $�d?�UM��Tz��P�<u(�6�b�֤� �e�wM�(��c�$��8r1{0>-j8�g'�	;�ɧ�Q�I�WQ�J��3cprQ4 ��+$'�Ve�2R}��H��y�$����t&��qշ���#g��޺Ӂ��_��X,�"�H�3J�����(�]dZ�6�'t����0w�L}�^:�4��e�"�{���g ����u4:Tx�� k&��J�} ����U*@E���Br�����a���g���!�1KI������H����`ϱn��>2�ɮ�\D[i.�l����٤$�~�@qܯ ��`��iG����� <}:wz�1EK�����:�K����!HRB�h�*V�2�A+\F�V"*iXi��V���+��L��_Tc�^���M�f�3X���g��x�k�G�n"��벽���~Y�q�߻=�bv���ض�zZ̳��*T�=d��Ղ�������'}��o`4 `Q.�(��[b�WF��� م$O���EL�c#���i�C�>��AW��ӕ$�w%jj��v@��y��\�EC/�����ѐ�6�G��%T(�9��_ц�D����.�m��sF���K�w���9V�8�mCnȯ�)r�B�b�p�{�
Δ<3�в�+?p�`�
�i%����h�w0x�?|Fǖ������:�>ڏ:ߕ7zM���
��"O�:������|$��2�$��?LN�C��hQ8鹈Z1�[0D��x��=c�lKQ%+�I2�8��ݒ���Jz��t��WS�x��#�YZLD���2q���+vZ�M��o��p�0��5,�f�)b�`5�����g�܄>d����t����4���a�U�W�g��ņ���j=���R�p'Bs�E�� �p����&'� �]��$b�U'}$��!��	�~Ot<��e��֓�M�/��Lڦn-�;�RK"��"g��/.OB��e]����
<�/���$i"C�J~㍌ ���ų�K�l��[YM��ؒ�$���f�$*1�b��A���F�����vb��/c�Fɯ̤.�sa��<��'K���[��2}���A��sۥ��g6'��Y-��c�GH����Y�}^�l��b��m(��V|�w	�[��MQa��*IR�E)Î�c�8�H��"�L�zx{�7��ح)&��Ah�݃^�y<rwr8t`"���l��o�J�*{�-1��Dp��g*� �tɚ�0N(s
�������Ɇ����L,@}dx?�/<7�ϳ�KY��n�H�ZU.+�e�A� mV�����Ԣ���x�D��k�q1C��1L�e>hR�t�?���Q�蠄E�{'���ȷ�D�m����>`��q�Lk������ѩ�j�5q�+�%H���JKw��a��Xq-ba����2z����"$v�	���a��9�%'��F�/9��P�)|e;�I�U�:�juK�5���Vϔ���0�p��5p����TL���!Xx�>���T�#��`ʞ}����_��Vh��H��C������!��ǭy2o�¶W�$D�����Ǳ\bWn�N�*Q��1k^l$�\;&�!�i���SpB"%;_ElO/� [��(�����;���d��	Y�W�8oA@�}b[l�ԁ�s�3�zB�����m�וϴ�|���/���A�Q�4����K����z�M����H,�W}T��n¸K��'�9�B#�o>�x��J��aI�Z��XG�K`��������dy'��<!a��s�9w�Z��p�����*����;E��P����#��
�x8����u�8�# f��;/}EW^��hv�U���mr���Q�L��U!�0b	=����qV���Z	��]�0Ӽ�Lh�������
9��}��0X��4����*��	�/ �N�y�{��F�\˹��|�tT���ў�&L�'�Cm)��b�������.�Bt���콻4��iyT�Rv���}^�;��Au�5a��r_�5G�L�TT*aM���L�Į�;�zԯ��s�RK|!���U6Rŉ�\H�N^����y�m��l��,ye�m�$�'�U,�v^��l�V�_�����K������TI��j�wc��įi��B�����ԍ��1�f�hRpN1��l�0�D��rr���	�h�Ķ{�u�Y�8�e`��wZ����;�4;�܍}��]<�=�C�����g#���M��Ĕ�8)���!`�ȟ�E0F���*�N�9㰍���  ��g���ky��!�l[�ۿC�EPCf
�1��pC�`�ծd�g⋷�A[z���
���x��t�n���ב?(31J�9���Za��o+�b�@�!碋ϑ#�$��g��:@�5�H �6�vx�ʵ����z�� �a��@�Uw���+�?$2��IیK���;���m}�h9��|����vr��,�J�Bn���]�  i�
��)L<�lKoΟ�wv����u�?���v��%^qӍW$�t�[ �TJ���.[X�&j{����r/����c�Ͼ�>���d���-��� ;1<��c�ӽНawA�4R��:��De�Q	�R��)F�39hl��O��K�C����i����j�;U��b�R}a��q�ڻ9ġD�y�]���ߗ��苎�FB��:���x?I �r�vuрF�/�œ&S�nF�Tbm=�4�S��ɪ��j@8c֦k�X�zl	ih�lRQ���b�c�~ͦ�l@��_�B!�����?�6�D�B�-��	a�Tm'�]"�C���Vg�N郒w�(:g���)�Z\����=U���������)%��{U���v_������+<~���3W��L,�u#ME��3��o����e�.N��'M5��+���{��:�����Z3c��Ciz�A���b��^������v�bm�����G�Kb� &��?����qS�-��
2�{�����\D���;��~��3^�;{���߇�r@�	B��i>�Zsvnؑ��D�O���(���V�̤�
��-w���7\�5�7��z����� ����X�вI�c�t۳�e�����:���&��{��}�*�;��E �޿���q�r�z�u�(�f=��o������������6�e��c{�[��c4��7�i��י̔���1d�9<��648�^L�p.D��Ίgd� ��T�(�w+���9���W��V��QrV&cʓ�^�9_6h����}v2�Դ�EJ[h�0~�{���>���]�� Vy��XDB[�����*,��[Z�v�@������zj��~x�o���I�H��OC�̬���G�L���aБ
�s�<�"|�;jVTe�I�!�N�͉�Q��VdF(+��St��+o�@�6%��q׺��a������T@�ۄ�6��n�����\���=.��rX���xIt����+r��7��U"��UHe���{��i�߃2��Œ�4��c��GC����3�j�8P����Q��D��w����=��3"���I�Կ�4�~��C��7\+x�;��$�� ���+?�R$����㽫�
�45�5�8~�y721>{�����6r��^TTxLF&>I/�-�G��\�%�L l<r��*r�,��X: ���Uj��22���ިP�:S���v%J�ϵs��_����"'+!#oD�]5$}d��_�!��0)�;�b�Fl�κU�����د#�f�}G���n#h̨>�?U��S!g�1Vqh짬�}�'Z��P�l[�q�i���V�˛Y5�sǌ8��@�=90�0 +N$8��g�:���	t�uC��WǱ1i�I�������%�)���r?�J��x!�\=�ߖ���W���{�@��:�5}��3�Ǳ���kU$�pt���yx� �@Pj�
�7�ɳ������ M�_��Q,w����Yǝ�}��P�����DX%�<�Q��#��h�B��ҋJO�cχ*�/�߿～s����Y(������y�V��eG�N��@ �#���7���*��g[�
 ����z|O &�?MYۓ��h�jg�^x#�z�Q���mp=45n�c}��d�?�C����Q�#�&6w�Rᠮqe!Ӭ�O��
!���+$A��B�É"��{����}9!"M�*E�_��6ɳAI$h��.���j߮�~�g�u@�٤S�m%8w��ݒ6�Y�&҉G��g�%�l��S�i��@��f���H�Yt�~[Cjy�L������DB� T�5�!���7��6��L��&�I�!�D���7�m6^&Z<tc��YpRD�qO�~��/�e�R)���"�r�c�m�im}1�*���X�d��?�^�""ǔR(ZS��2z_��	�!tm.��d�1���z�1Ư��
u�M{�Rp����1pl�M�/Y[F����T��)Q��U���׾[�@@�M>�4ײ��݌��Oxs/s(�Tp��	��l4�� � ��l�ױ�Y�|z�B�1_�9��m�� ��&;N�܌��x?�҄�s�.{��Rm#c}z'yŦ�S@6ҷ^��P��9:����Sw�^3���kW���}����<�� �f �]���0���?6Wjy��\8��j�Cm�ڍ;��\b�g����� �S����[�[�A<a�׻�m3I	��F�*#s���n�K���X��AG��ƅ���.�I4�7��h(Ot���q�SWS�Sbh�an.���J;�eb:�L��"� 
�C6ע����#:��K����r�Zu�~I,�;A(�������{����h�aO�+�>��%��5H�f�(ь����3��$>�١�m4i(�mծ��d�����n�c�p4��-$ku��+�c�u��Ioup��Gt��x����7��{و�+�����gW��Ɣ&�9Ĺ��\L��!_��1���dL����f���1�0�[�C�}	�F��P噐�	����F�(�+AQ��*)o!����3��[�]{�ErC���R�x��i.�+�j�iZ�^���$���O��-c`d�AG�5Y������%�i��UF������1&�����{�5~v��#V�ՑĢFb��{��<��I�_Z�u�n�6�D�M�ol8��?��WI��l��a+�!�	̊K+�#�s��N�H4K�5�� ���z�|�|�t]i�~<%�a��L\�
r�����0΂�Q8f?#
f�Q��4}�B����I"�~����=p�qױ�b	l��K�@�88m�,�`;V뻣评j���n&�Y�F(#I`��.�t��Np��Juh.�C�m�[�mX���ň�rO���
��$7P��l�;Nf<Oe������ku�XjyT�+�3��aT�C�.^)/�C�{taS��H|��$*g�� ��~�)ʏ{~�j'50�]ct7����������:�:t�H�M��7�Gq���3�}:��r��S5�`�9�D���p}v5�����9�=�*��L+m�P�aE�M�P�) �܃"��
�/K�t�>��I�v�gP��7����hG9A�T՜���W2O/�;��F!)Eh��a0�����ܣ��<xd��%�7�{��C�Bٟ��i�A%7v��"q�k��	��O?S��`�	C�ԕ��d%A|�^�s"��n�=Զ���}8Mz��o�������޲�Z�dw�a�O93�T�L��Ν�!kq侮��[ǽ��E�w䭋u�p��|�-�S�t�5���;-�R���sw+;�L�9lG#�8���l�\hF����EZ:e��ig�?Yj�+�&�������Md:	�)4 �O}{*ykbE�np@I�{p]P boKckMe5@0� �띦n`4ǯ�h_�w`(^<�Q8K9�?���/��J�;��.�&�§R�R�w�%�(e������3?Q�	�ה�u�������1q�6B��<#�>T�1��[�|TZk�������o�AݖY�-5p��C㗡��J�Ny�?��)���
q����`e��u��7�Ě'�4d-R��v�����v��_π�r�����q��:����9CLk�9� M���j=3���r�^�f�}��݌R-rЖ�¿N�np	r���	eҬ�֚�l�����E-ٟ�EL+7��l�;�^G{z��wj�à,�_�O}��7�jn���1����R{�I�>��/ �溌�Eyl6�o�#��hL��"/-�,"c�>�734�7��rfZ%�S���,�*�[��xO&ٚ���\;5�½�W�eT� ��=�#����<ɣq\N�/���0B�FK*�� ��$ �}��QB|@���D\�z�#�L�VEC��mY�]|[�`����9��%b����G���B�z��)��F�����!Oќ 9�Tt� S1��p`�D�{���ZcV�2��nkiJ&����\������Vd�q���e��T2W��Z��U@���@�Z� 3'� ��4���f��ޥ��ep{����T��KșJ*x1�ՐrQ��	��M��Mi��nv��{Ke�k	�i�o�pk#q���W�p?��spV�z|X�̌���h��|��2I4���3��!T-��t��9��R���Q�")�Th�ܜO�ge��? ID���5Y�;�,N�k��qd�ɨb���В\~K ����
�<��Poϵ�7Ө���V� ����zߴ�L���z]%)�BGF�(^��F��uf�&
1��h���G�2���ǜ-O�pj�CK��Sgڽ���;�����B!Y�p�����[����sI(���������e�����o��@�cw������W��s����5��@�3�9�������
d��!��>�+�# �W$ʚ���7�_�%���<�Ϋ��j7����(_�.�@\���16�X�sZ?8`Ȍ���3��U�%�r}K�4�ix��P�CP,g{=CQ��Rk}XuU�cJ@P�PK�Xfւʷ������N*7TH�s��+Š���ף}&tj�e~S̢��&_���Jw�O�N'��j�ʵ�qר�uN��3I�a��f��L0Z�ækl�ž�j�"�/����T�\A*P��B��U�fc���\�v�;V�����TT��Զ�-ĥ�/_*I`�ac��Qy�9�OR�O�q�;G�k=I�GL�<'���9��۬���L�&�?w�x�v#��.�i�옴,Ӻ�j�7���S�=����N��.��qtf|�og^�[����ư���疥��ɝ��Z�:172�����7����m�]���@�<P=?�Υ�D*��t�:�.]��۸��*\�V�˒qd�ɟWɎEÖ�D�E��Ūv5Z��.����9�*-J�7����٥����/���N QVw��u�ѻg�/�1ɇ\�a��]X��l��Ȥv|�N?�1iq]�:y3���������,[4^�p�?���:m\qj���e���5`�2*ph$g�PWp�|�HcC��2�6��.s+�}�D�Hm�͗��z@����r�uf'�| �Ƙ���(!މ�ݛ�`Ե�2��G�i~oK��ۋ^�̀�ۋ�b{���J�u�1�m���`ŋ�Gs�x?cY�ߟDKz�z��DL]�ih_���8ߣ|:�~ʮ�i�OvSJ�+^q�h%�'_�I�@aA���a���8mw��|���rT�՗/a��y2���B������ Utl�rɌ����ES��Ĵ	�m������,�����B+K���j�,_�3#�h�	l�w�s���9I��j�5_���f!�F�B�.��ߐ
B��K�+�?��,u�*84RV�.��pY��O��k�q}�! �%�A��hȴ��9�/S&͝f�j@�2�Y�$�ھP�L�����A��j� y�������S�������g .9�b/��JE��,��O���O`��Ɛ�Qh��%@u[�0�=�"�t��6��Q�	~G/���Ȥ����5F�)�ڝj��-����#��}�)	9>U��U�H��W��l`�1���u�0�]pA�.-0�C$7������\��t�1�Ad���z�Q��5���0�| ��������00�O�a�*�B�5B`��<���d	���Z�uC�n��e�H>������=8,�KWH�\�om��7?��]������w���ꫲBy�j��l�� ��Z^��.b����*r�)z9��)5����N�a�N��h�\W��@[�AH��ş�����`��G��?�!��N��a�'������S�w�Fs#��H�~�h
q#�n�ӫ���r��W�^A�CoM6Qo~�{�2 �ݑm�P��ǒ���=8[~�i(Kh�_���Bl_�&K�}_��1���m�
$+�Q�d*x'�P�֧��n���ZǓe���]��N&|M�"p���_�_�;I=sX�z��|�5�e�����̶�	������M\���8��sQO6�^���;��!/�Y=6��Cl���J����]�s����WR��g�=�����R ��?�:Y����	��k"�,�����P�t~B����@�Aٟ���"�k}�푀,�>L�^pE�C���H�����`�m�}90�4�T������!?�[k������y��1{gc����~�r*9�ìEj_�45A���y(�2Pt�"�iIZA��~��h"��G)Uq�|Y�����M���m�Av�)���sG��c����w��w�uMC{ߣY=B,� �Z29�)x��%�'@(�m�3n�N-����_���AO��0����P8A��EgO���KYC�n��
���4�T�2�P0���<T��`ξ���HAg3�?,�@^ķ�����s
 W���OUi|���ih���ΥZ`7�+�7�o��ʷ��@�b&𢠄��Lf���8��,���m*$u#��c|Ÿߪ]�AK��g����sW�1~���L��*`�CTJD�D��b�*\yE�Պ*6��Д����n߈��%&�Oli����3�4��q�����\�u�A`��i�΋hI����;�V�̧�#u�z󏢜]@�Y2�M<4�x���a�!�~ip �m�O�]k=ki�oS�mB&��A�̞|�_F�n!��Ñ��}�V�
�>/aR�R�|��ah?sNqv��5d�]Җ`~+�⧇l�j�<�V��RvU:J��jt�4*6|G��Ul
#t�y���܌��H���{T?2oDb�܆�=aN�ܐ� �������sO�֐!�����J�2��������4~l�fC����>�2�[#'���L8�$��pa��X뾃X��7�;����8�z����i��DK�����]���rB��|��d��E�����Ζ��������Sf�����������W'�[y�ua&΢���iN�RX�	f��w��g4un��'��߂�)�%�ۂ����Wx����F�T	��C�NƲ�2�f�x��yM�@n�8�M��ߦJj�Ђ���"���wژ��n�%̃[B� )��^A��)G���d���P�	*5����������k�f������T�&�;�Tl�'��l)�ҎȻ/�Ͻ�
?� F�d����Jy�&�g\;�1?O��z�m�����0ENO��{0軂6����Jw��t���:g�� t&�߽�H<�l!�}$���
V �W�B)D���@r������uZ�0w)���Vy�� ��̸x
�[aO�c�t�K����4u9�)�Q��ޮ�� $ׇ��6��{kb�2g@x�'6J\��D|}[уxM |y���+"�^zyK��c'����Llq�-��v���س:w��:V���)�w���,�U���5�c	8�HP���,<Ǧ�Κ��j}0��j�d؍���4� w=A)�y�ɜ#�xD�Vq�� �z�Ɩ�ߑ�v�&̄Ƚ�q���;1ǽ�Ȣ?�����۱+X^U���썽/*�S���ߞ���#�d�����,���ւ�<������tOС����o`��0�������RCИ����"p�G6!yi���	W�M�B[A56�����=���5���w��8�r�m�!1l��d��Q��32`ɦ\��l�e�U�M�R��m�c
��^�g�ޘ���)��.xgp:����J�/�����SE�<LX�`>�ԫ�{7>:�)d�ÚnA]Uj��`�l�j���������!p`@&�!{�w�ܾ|U:���� |�t�(�x����N�$��m�+Rl�-��
�>�F߿zL������Գ��`֢�4�� �=am��f �c+�o��b�py7�����u�x�ɶ�nj�Ok!�>���4�ǰ�'KX�	-휦�ϩj��4N����u���Dy��@����m���6�R���F�wE��7��sD-̞:���qm(�P�͇����1|lZ��(��q�eO�!��%�Τ��r$��~��6���!{IF�^�#�4гn�h؋���w�b��Rc����U���^����O�{�("~&�����ڄ��:�#WR��do����K�";��>	G�c�J}p�G[h?��r'��}��{=���ÄK��gN��_�񘨢"�e���e)����YQ��D��W�큃���|'�d4g�7Pq�,�>���X�*H�wl�s�-����x�:"(��ՙ��ԁҥG6F��/���~��C���.m�w�K��i_^y�C�5�Ł
4���Ưz�F�!�)��U�]ʔvv�3�K��J�b��H(�b_\��W�z:�T��Z�EYZZ�zr�j�{��9x죃hPݴ�� O��ξ</ȁ3��j1��"��T�^��������X�n�w�/��	?�5��"#�3��MVz�8>��;����޶8F���w6g��k�cE�|�R Ʒ�->yCD.���$��K�L9/~�ϙ�y(��F(	ae�:(�$�.=���o�x�aа�S���VT{E)3��b,���,M�W}$K����Vd!�x�`;M����Ur�ؒ�d��1�O�Sӥ�rK�fQ��1��.Fw�����-v�k|j�k6���� tL.�8��E�K���}�Y���k�ړ�䒭���5@S��4�u�����x}��o,��P�8�^?M`�~�ۅWr�u����ȆP/�B�(�r7�}�0n4<�j^(��H�9\)��0�����Z馨����?�e����3�l�P��Ðy?׾�O��$ݦ¯���[9�onU���������y��8D[ؼ^0�2�{]���\]�T1�0�M�C 8+��E�k�5�ϰ�Ʊ���־�8&G��Ww'qx���J$�ul=���ʬ��!-0����g�hڿ��3(�^�g�).#ڢ8����%X�>/�fB���\< &����mr��'�����jn�֎
���-�"x���g�uM�H���Ud�ϵ;H����o����vT�!��%P�	��GtY�+�T�!�*N��$��N�R�g�����U/L�h���Ԁ�_Y8|�+@Xj��qYQ��l��[���{5߹G>.) ��\:��ƳV��t��kWh��;�� g(��L��y���?"�B&&n|9.MB��D1 ҆��sIV���؝�YLͽ��f共����U��,i�Ĵ�#p��2ng}��(+��e�I}�X)��yx��aK	�+352�ϬL�O����*D[�sSБt���ٿ�2\��� ?�9��/���)SXU�k��#Ff:g!Q��=eٕe1#5;��[�_�0g|��T��sh��@Q)���e��E�=� �9�q^I,!�~��.�Q�<��������W65�*���BJ��ؤ��sv��`�u��y�� �>���&%�e��$j��w��p�8�PDP������~��1�YaEˡ�hd����촇߬� NҦ��������� �7��č�#���Y�7��d�񹎐x�E0T2�Mgm�?o� B9��EϨGD�y���������7�75���^���|�_ha�oa����{	i�P@#XZ�e�8@)_gٕ�~�����K+�a�mC�G��%�Nu�E�Bȯܦ�S�pf$�Z�d<�� ��$�j���R|U翂xS����ʮ����u��&��8'��5ʞj�b0w�0��W�%�I�k+�����</������V�xa�Ξ��b"���g�O��`��)��_�4.q�~h��^G��\�vu���g���ɵ�HX�1Y?�Ʒ�c�.;}�SN��&�(<��2t�J�+��p!*b!V�0��2��V ��lR�(��"%=�4z�]��qO/5�Tn��VU�F��p�����k'������h�n�<y�e�a*���tq�5���J^��X�M�ݗ�I_��ė��=�������V��ڰ p߯����~g,�bG0��*�ks����w�0M�;\����!�m���!�4+L�_�1ť���^�>0�����p�r'�G!0��_�p�6����J�VRL*�l�G���Q�.�	+����f�P���X��ȐO9�J��.����R��[���_8�Բ�ዲL/P��T8���#��Q�cUʣ%��\L�M$3����+���T��W�ՆxĂn�hr���tЉ�{��:1�	��zv�<�r�N�9*�6؊a�0n#�^r�P�L���-���	
�
��;XS��KBP*�b1���U^k{7��O��[�%��B�@�x� j&Ƣ^�	7��k�1�ڼa�M��	=���J����A�Z�J3��I�8$���dUÀ��i�S8֒0�o��:�j`�91�Y��ǚ���y"Mc��7W��F�A�y]����>&	/�(�<�O���]�0�b��5�H�i�->_ܢ�s`U��Z��CI!\��#R[M��g�L��� i;��I�%w�#���	!��4�%��}�oMA(�c辶�S�w*ƌǡq�H��Q��C  6QX,@�(�I���4��3>ƍu
�Z��`ma��B�	�5���)�^����~9��K1�%��ꓖ	�pr4�-Nm�t?lp��bO�p3��Øc˝;*�,�_�44����0P��R�9>_]�--6��=��r��6����!2q�di=>����5�g+�IW��6|�©�"��bon��&<T����@U:�K�|G�ttc��8T:�P#�H��a�^Ԝ��٭aV��垝c^�4�
��/��-�d�j�a�~������q/�<�b�Kf��������W���EDK�X��w�M8��oa��幛���s��b)P�� �s�����B?��R"�E�t\�5���XFx�b���M���2�WX���I|XB��@�S���^�Wb�g���Z�����`�[M�ao��s0�F�։��"_�ͪ���6:�(��(�7CUz�����#w���Uf�|7+��h��0-�u�������_�
P7TP�if�đ9Fl���c�㥣m3��2S3�#"8�0z��X�&I�Yw�F��O�~]HP���u�,�G�S�ʋX��9�9B4J_@��D/)���6V�܁+��>~���v�4;Ȕ����JÚ�}����Q�Hq]� ��X���]���ka�{�:7�Y�V�y����`��#�}�K�HO9��<��`]���s]���:��%�#�մR��ůT0���ђ���](�$�ƞ�����x��Yռٝ�������f���Si�Y4���� t�_z�lE|Z�E°�V<:Y��l�p�g-�}�B��1�#��9�G%%�p�������qܛB�J6�vu8%��|;��{d�=���6Hk�>�x��f����������΂��)-��K��Z��8�'_|V,`���D���Ի�ꂈKw��s���ٖ�vd���� .3f���~yۯ�-ay}����Z��%�e��y2d�@bۊ�yd-�b�zOϜu��� ��L'�ʌ��@j�@��t� �����~�~���6d�_�"ɛ���{bH���^.Dw��v�c�t�FN<��Ȁ�ە�V:�.�?d�t���1m�#�	 ���
��3�U�a W"3}�"�F+SR\x�z����^3|-�/�X���vzG?���.js��naV+���o���^}"gO �+ r6]�����#ES�7��K������lU���]A�0AȆ��^P�5�*��[��%��c�
W�cimn����GvV���SBٲ8&u��ĕ�Ӛ���%��T+��n�]$m�r�n�Sq��8��+�!+�m�9h`i`����Ru�H�אּ�*B2P�a�w�d�lSE��`����$Hʝ�Xz���PW���Oq.d��W��/��H?��JR#��A~�����sЩ�����;�4���>w���P�m�ȂL�ߪj�R��r4�w�`Q� �B�(i3��z��V��K雸>��>����7��ja
�IEq���������R�����/���y$WR�-��(�#"�w�^zt����ی��%Ta���<:��a� 8���c��d\�"��RL��U����h�/#GFtxWbS�����.CY|I�2��p�E���f^-=� [�"��u��Ji�t'V�-HڨC�-̜��)T�:~�L��}���W����w�-e��u��Y�G:�,}������Ey����/pb �?~:�"�7Q�0�z0��;��?Ê�( �H�ԁ]P@��?V�>�˕!�(��aهy�����H{��{U��Q��ْ4�|e�Nޚ
�fn(5�����9$��)e;�Y3�#CeN#j&�o� ��x�T�- �<ÆR�8���,%�
���3b@�%�q0�w**�������_<~$��]�[7m�x��d���7FN[�lVB�&��z?N@^�#ط%33mGZ[�ב�9ؕ�]���"�Tƣ�~)O�4��]�/�h� i�_�-R�ew1�:ݽ��|U�zש�4�L�N1��8���݁Fӂ'��}���^�t)�8O_є:T�(F����ҶT����,p�����(�{(��Y���Ԅ�� �C}X08dA���u�6_������������Fw�����$V����/���9�%�)5,bȂt��̱/��FX�b������n���������l!Ղ��X��9��u���� ���,��Q����*:�Ե��YeٴHK6{!͙~jgٟ��>�nG���M?�m��p��Y�����U&���v?{�_��D��ſK����=2zdw��&�x���Q[�{�g�|kxk�ĝ��UI�tm��g;Sj�Ρ�Pi�y��e���C=F��}��j0բ-x�Ɖqb�-Ab�["����<Z�!��pF�R�Erp-.���g���K#�����$�i����&��ww�?v��n��vU
����{��3����y��_�X8�o�*�'��Ͻ��K������}a�L~|��Z�]�?|$��
?��MX_`�r6+�)l�E%�K|Ȫ.w�q��ɜt"[�ĥ�d�z�q�v����t�G��X,�'ɬ���ZW�T�_uwg	V��b8���Co��)�y����@~� Z@+b��8E�x��e�.8v��Dv�=��$�q��B+鸃)��ح%���~2U�/��q�������QΦ�l����nsUfV����־/u@�X4���;�7 0��_�2��we�� �_CEh�g���F=�oN�I��<CϞr�����_�~��J���"Z���Ŏ��?��&��:8@��ԫ-�i�' �z+5��+vQ> *}�/Mw�ܶN�O�n�]�9�������ӭ4!��u�𷇮�����1I]I��J�&�C�s��MD�:�.��A�S����h[���l�~�ɧ�P	�?�5H@*K%���ʣt������֔sT�[��1àe�D
���2��&��IN�v�&��Y���fP`/�#b��X�%�I~l��O�Cr���f�t��N��� ��g77Mp�����4����,���{������ux7P{y`��fm�4�}<.�!Ѫ�q;�i�D���c��zj�E8�0$]o
N���y���_�ctmm��hȓ�&�R�2�)��Ÿ�/SE[-��#ה���*�T�YQ��WA�����
o�M�ԡf?̵�A��o�j;�uG���5}���d�PWKam7��H�u��TDa�\욍n1���`۞��ҟ/: �z�����+�fʵ',#Ee�{�o�9�]�w�ӯ������/a@[9�VYt��� ����y����D�>����
���	�+n�$����bm�ਦ�A�����Bk�.{¹��p6o3�ڼ�;����	����B갆��s�&�h�_�����H���I�M�j���>㺪#�B��,ZQP#󚿦c_��x)�PF�����2�����9(�sqd��e��7�d��ٕ?s_�wA�fțo�`ź03ӁA�	Us:y�؋�q�WG)CӈS�n����=�f�ߙ7���zZXbS�}��(���p�<�B/�;�Yl��{Md)
�Q{�h���Vg�!z~n�b`) ��v�}��z.z���5E�c�Li�bZ�`�'�e��j�⟄����?�o(K:ļ��#�pk�l�!�x=���W�����5j��.0�I&��C7	��7�	Cm9���Q5o_�n�?%�굧'�e%�M'��9����fd�IO�k�f?rx���!����;��&0�e�$���]H�Es�!<�]� �����m��퍕Hy%���j�A��me�e�eM��w��H�t�%�5�eCS�����1�p��YC��'���򬙁\�"%iUS�6��a���
,�H�
d����ne�RUx��$(T�[[(�旲o! �4L�M����N�CBYj6�SB��/X�#��ht�ix���T���tZ$6���s�tR���]��iP��q }�D����[���x�����˃o�������|� E�|���շ^��h�a�V�m�J�}�hN�����6[��!����ʐc��)#֬`��׳���D��ٜ���".f,Sf�F�)��/3q�{�9�l�+z�o*�m���H�j/s�Y�/I�Q?�I�vg���<�5B!���?���L��a��J�h )�1CGg�K/����G&�'�)5Lb��aAzS0��)��~��z�Q/]����T���'�>�[<��"��R#�s:\�яŠ�嬲�g��/
�^G�1���&�d��?7Qz_H���#B�~'[d�0�Y[C�ϫ֥ZgiK�ג�Kt��籜��`O���o]K�����ƔyS��zb��͜%�NAW��3�%��ɓٶ���+[xY�}z*.����n�������.��^<�3����Q'Mڠ-������"�OG�ü?��X�.a�u�����Ƈ9Y;[�BD\Y�?��Do7�8�-�"r�ϧ�ed�WǲJ�נ�0���%-ِ���m�V���0���4J�xEnFA���\Z�N�h����@�
e슰&$�ѱ� " �|�� FY�B}zY�n(v?��*X�v5|�05��n�{��	��r�M��G=7)ne��)���)Ob����ʤ����5.A��.��ek ~f#�E^o~�t!^��hc;��ȇ��d��E�Ҵ`�fgP�gTeH�%S�xi��SԼ��˻<�� �F��ʅ����C���i�a�X� �=�/�N@���#�b^����*��(�t ߘK�M�u����C���̫����N�,�5B�83�~W�����f����r�܏Z�7�߇�sq����f\�Ha��B/���G��%��*j>��>ma�����}\2������[w6ay�#VA���z=JJ�A8zR
y�B�W�Uz�3tڒ{,�G��0U����Jkk���m[��F�&�V���S����L���)�L>�W:���~!h��דPc3Lx2�1@♋�L3�R�)�e�%�{NN�ĒC���}Y}���{^j��ւ�))Je����n�`��aF|+��5D+׽Li-��t�\���F���\5w��9@�7��Yq�QM�+c{}��W-�1��Z�ݙ���%��![�D]�ek|���߿���X������ӓm���ƿ)���~��˙�SQ���d"Eݨ����l��[�0����o� �3���.�s�:�aj�����{Z�G���%�?x?�N5�HA����`:�.�\,�f�B
=�'�I,�@�Gc�2}�������pֲ6�H�����ڑ�i1��|!Ur{�
u��
����Jf�dLdS�NG�hyd��$)!.�8�����J�¨��-��ț¿���̺X�׆��wc8Db2w�t�y��~ �9Q���e��Cf���>Lۨ�D���c�4z��X���b \)�fs�C|��w�P�xc��e��q��҃�羹�P!r�o3f�Ӂ�������j��Qg�P�� ֪�2^���e���ߝ*{��6KP��w�AԺ��g6_�l�էK ���T�N_jY;��+1M˘����}��K������#E��=^�OK	י���oD��i�	��.�-;E�rbu+��5X����-4�+�H��G�[p�
�_�41�T4�tW��4%�<���~UB44�������6���ү�F6
�m+:r�w�|��2�l�R�3�V�/��4�|`���庼tJìW[����yp�q����F�x����=D.I�+�_Uk�#0�i�A�Tğwi1.�����^P��CaNԗy��U�ʗ|�v�|�*�F�b�-��y��#��&�q�b���n ����b�b��3-�I�,0��_���CA�{J�<|]tvs2S���c�^�����W= �:���|`/n5A\�]��ҤL��4\�V��l�R�Q)5� �=���ܘDO0K|�ɇɋ�U�Y�;d�Ә�����~�`"z���p rk��T3�ě�S�cA���D�KO�x���Y�˴{6�q/=�`��ڝ,&.w�!�v�O�Q� <s��]�o��!�՗��۲i�#�~:0Ї�+��E�XW9Lr�$�R��'��$`w��i��������e���u��,�y�����T�@j��\�O%����O�r�f#�}�*�o���{$xo:��Av���A�y}�����.���sQ$�oD/��J�?�ڦe����_U����.�������)/W�������T��D���"���h�Bǩg8��un�-q?�72����/ȑE��񫫸#���F�&��ώ�^��4a�����5�Q�sȎ}��F�-j��+�3;L%s���f^[0��D��+���&�V��`4���y��@@kPW�*���]�O�.�*�Q�+ZR��q�v��������*o��څ�1p��T�p�t�=�B�;����i�[M6�ɳx_?|��/���c�+�:�����y0�qy��d�H�k��>�ݞ����`{F��m��p���/;I�9uh���-hm�'t6(R�DI�/�'���V�J�]�Y���J������4Bg�EQH�(csi('��'h��^��DX��{����>�-lw��V�P�	7�% o�:w���P_���9�Eg:
*z�����W��a�Nt ��Y��Zh��I����_�e8l1��K��*3���^��V��t^}�_�Al�2�q�P�q�Π��a�/��j����XlA{�dxuۑ�n�Q,e�Nf�X����ЦE_�?,��h ��c�p�9�=󴭢���ԅ�g0�sO��<?�5�)���d6X��*I~�B���-�����4�.#�K���[&�G��=���yо��8��T�80�م�}�#6�n�-f�E��d�!��u0�G�ÿzk��R �S�?��Cw���ڗ<�{�I�k�b|���z����+��_D��D E�d�~�v�s��������<����w_[rG��oZ��f�~ �
���6���������X*��W�([�K��iP�(t�)��5�C���Z�n��ˆvE~"
&q�~��s
Z�ß2�Z�3nI���)��i�%�b5�T�ap���%��=�x�v�g�š%��~�7[�]Ӑu3���T�<���# 	�L{����>�2-��0a�V�>��^���un�4���tK�<d�j^���j����O�h�J���FG;#���4�Zi�=q�P��hX�/5���Ȃ��3܀D�=Hh�[�g�=���Ԥ��!�����i��#Ͽ�U��ܔk�\e>�f{�If�a^�X{m�y��W���"��qSwpý��Shf������k0��i�]��ú'*=�]O�e���n�m����	\K�JN)��1�G]`�pm��� �l*?4�-��2��q����N�����cU,�niH
9p�?KcԇN3Y.ɒ
1AIq����8�稃\9��i:�to2��MK|dYhF��S��7lў(y�� rJ�3����g1^�/�Nh%WV�l�v2�H�~ǆ����`�$��O�nA���.��a�)�B�� h��#������� M���g�8������Z�$��$a��F���(T����!�2Ms������3�l
��N�ގI�P`�T���n8�}��pkF���RQɭ�!3�Ȭ����?Y����3I��9�����]���t��T�M~p�c�r^�:�F�v�FU�]ǎ�Z_{*�{[8�{`��3$|�5����{>V��|	M�j��C
�1�i�ކu298�Q�Z�B3h1��'$��3�ً@S[�|��;#fU�����A�yO��eq	
u�V�fHqG����K�y���r\)�Rt����$/lI=|-ٛN͖�)N��-�w����/	i�4�9�Q���q��KO'yLr ��e�MNx�v�0��eA�N7�l�B���z�ELGݤX,�sk��p��>�[�JOy�!(vЭ��/T^rz�~���N��)wuy�DL�H���J�0��M�Lg#mh�� ��F(���� �{��t�y��L�X���m���S�)��U07�L1K�z1C��,n�.�s�og�Co^i\��<��C���~��+7�|\�bNA��]jI���A�B_J�K��=v��`��7��*���PKgSw&߄�CQQ|i�4��l�R�PF!��h�J�R���:��-Q'��3� �Û�˂i��:�[�Y>���>v�C�#��8FIM��֞�{A���X�l��6�Ӟ\LH~$���"��Rf���r���WՄ��T�HB}�p� Q5eK*��$�X� �7���W��Ns���(��~#o ��ڞ��t� '��4�^��>٧խ��$�[�+Ϛcd�C�\|���`2R��<�-�� P���b:�`R����T�`�����dz�v�|h��������F"�Sm��NYF?��''[�`�rcPr��}�f#������	.��cݶ�B+쑄�;��=:�PߧԹ��2���/>- �lI[T7Bt�[��2i.gH��������=��Ϊ���?�Lk�}�*������A>8G#�A����2u��o�X�5u���j��n��w4%�A�E����6}?&a�s�ca'М6l
7{ ݯr��2@��֧M�}!@�w�)|�HR(�(5Y���J���AQ��6��KˊL�_�F[�m��B�T�̋��YNIcIn|��a�t��Q̵̀i%Jp�mzvS�����Mq�Y�h��=� [ !Q�V�o:@.���ˆ�p��j=~/Ⱥ�����9M_o.�w}=��^G�3��GJ�y�KU���J����N|Rf���̰2��x��|�LF$|��U�q���)���ފD�Љx�0�N�2�3"�.ÆS��`NCdY͒[�1M/m�G�/)��9~��^��.�6�v4p����_��-x'-�;�<I��x��B��Yw�U�ݕv�į����Rͯh�D+�vҬ$���S�WbB�-�|����P&�q�t�@���2�*js��T�fĥd_�=F�g��X�Z��5ß�c��f
$Um��.�{����q2�;d�(!B����uڼ��坾R� �<�yl��,g�*���:���.֤Q�oC\�C�s�)I\T��8���&�+kU�7yVBE�᧏��Ep�7%�MTxF��M�V�{D�X�
����䵑��̜E���r�a����������^�.�ɕ���j�JW�Mv���d͸H�؍['�)V��Gc�O�1�H�`� ESz)c�m�@�d�NOm���X%87˂�� �lya�	�CY<�#J��gy�G�9���JUa��qȥ��|�W��kN��M�(�������d��.!��H�3��G��)�I5�����ūp�5X�w��z缑��,�,Y���1�بĿBi������l�!�׃6F��yn=�DXCQ����8PK���5�,�8p����kp݈��@[��>��|����0����='=�֔��Y�*�m|ׯj�L����3�٢�6�<lN7w����9��LE���8F~���E�
s�EWv�@�柂�� "P��G��8������Ǌ�a��a`���3=���iMʚm�M4�KzdQ�s�I^ �t��#��?���>nR��'	0�|����eB�� N7�zB󲳽"#����:�¯�T��n���ˋcr:����b@g�.ˋ�C�5r�������;�b�r�g��>���xi�oϦ��x�R��آ$��9����O,�G����y��g��q��=I2�9[*1/Wz!��,9S'�tn�>��_NL08�<�ZM'i'��UI��n{�<�hN���\��N��|,�S�P��LOI�E=��*]���O+Y�d�+,�R�7���)��S��,�$���S�*�:��K[�𭖘Oޭ)V��4f��G��;k�C��p}�dޞ�#�8�P
6\E���f�]*1ʠ�u����G�C�1<[��x�^�����w�d�S�c/73pW5�K�� 'PX�ϓbJ�_ty��FڴĮ*n"�e�4W�&��Z����^��N��_�ZXB�J�yCS׶�/Ckfxp��Ѧ�b���q'�B�Y,`m`:�6�n�q�Y�:W̪N���wN��ū�d���d��8@���G`(�Dl��0}G�n\@�6����[����U��y��<5>��aJ���ѸT��9\=��SF�A��i��ן�����t����6�c�_bPzk�^ͭ2�'�~�6[������%�G�c��tAB=�R�v�bb���v�ͥ"C#yZ����ξ�X�q>1!ϋ��>7��΢*���K �~��|lv�]��<7��?�]��a�0�'I�6�C�T�����Q#D�f5���s�P��IJOu��LZ�s�d �g�0�rʰ6k���ڄ\MiJ(�I y�>)bk;�͟��0bR��8�C+��H��]�G;t:�S�+oY?n��r�Hkt@�먂GT��z�RwmvC��Q���90@4��nͦ9�p��?gp�j��.�*V�w�И؁���f�N�ǅ��BH�X1����@���8���ƥ�v�6}Z�G{r�s"1�B�¦���94<�ug3J�����M	���_���� )�a�v6�Q��\����}j�_B=�&���p�!N>�CI�9�X3�+���\kD^���q�ԁ���)��e������A`Z�Em�QD�ofT�'}���Be�d:m�oq~c�k� X��-JR@h3>�5��Q���r�����̑��:@�k��\�1�C`z��%�L_1{+�� U阥w�R�P�L#a*_kmb�����6|Y�'؝I��NQe�؀��L���u=L+��m�!j���XxSU>Wx#�y�ZU�:�4���̑�����C�I��
I�8�u���l�a�A��T�$��j�5�||�[X�;�3u���Nf�˪Ϲ���R���R���.f�!�G~����VyM�t��h�:��k�TW���G��_�2� jD��_��u��V�HLފM��!?0�J7?�i���������j�1������20�d"��Wn>W�NM�r\1t����"�I)����gbH���"�U�3������8:�_��rg@8�KǇ��P�@��Z�������� &+�z��͖[P��Pi���D;Ƙ�7|�|m�?����e���Ӥ��d�뒦l(5��"N�:�I�i@�_�2]������(�NF-���d�)@�vj<LD+0�U��0b2V9�p�co=)�iy3v r��x���e�r�K�vo�i��_�Um� J='6�2�Nx�>��#�<�ʟ����k,�R���\'�y���b�!Г 4�M][{����Z��IQA0��x��R��([sZ�t���}E<�{�#�Fp/�j�Xy�[�{�&X?#@��PH&�D�Hw�My�u	ֵ]��N+S���&�<K�U�k;GE5�6ɛq�)���w����!$�6��tԌ7��%\>\x*4��>\п�a����ꦴ�����_��
AJL1L���?��^�(Dv��g9�J��6ͥ8��,��x��=mu#�p[@�^g�o-{���{�uCa!oٱ,)et�l[��*8��z����4K�17�G��l�y�Ęt�`ығ}f�5�;��b&�H�Gh'xS5vj��V
+hn"3q��Q�mn4�ᡊ0�v,�ө�I�t�x�넺�$Exj#8�Rp��A׿���������~&��kzn�E@=W�k�>�(��-M�LU⭫I�0䅤�=�슧]�J��5䷀�??��gmͶv���NX��ג�<R��y+f���Y�4�մ��$`oml��ї�8
2sh�Y��*�٤bx��C��í�Jh%��5٘\�x��ȱ(�x%��柵0ϱVc�Q��ռe"]CZ���׃\��T..�!sVԚ���
�U*��rv �\I��>ˠ�J5t�<�`��yD����c�@�^N�VMU+�{��.uE��D Ȱ	�����u���Ԃ�g������X���;���v���"׋!�J?'� n%�B���Y��N>&���~�S���^ T�,�������u;������I�*��s⥀A�tA��=�[���'ϫ|�_�ۺw�&EX�p^���Ӌ�qV�K�Kj�:���J�ka��9�*��g�NF���AIw���/��L�>Y˙^c�t-���-J�%T(V)V0r3���N=8FCZ��
c3�/Ŧ�g
X�J�h�5�	j�7A�YH��q�wꈞ���T�-r�>	���[�*`$�J��Գ���)�yO� ��/4��^�{@�$~��t�iQ�q��9?eezy��@@��r�^ �/G���~�n�U޻�!5��ܹX J{�W�5`ȸv�Us�/:�Z�M
T�}F�~4. �B$t����Kcf���ӭ����Cl��wX�C�{.{ҮQp�[4�c~U�X��/B��I�?��0+��u~���6f��/>'�H2Af���+'Ah��|�J�+�?'�p��PJ�z������#����w�Z��g���y?�)�g�6;�'���Y�+��U��"�� �5fOڕ��5�|��a<`��>T`
[��m��Eu�Xk��	��0%��*?��Z�8Ч�1}ѵ�MxQ��\��{�Y�M��q�V���Xs]u�O˟�:`8*��a�+���/�<U�l�����F�?���� �d�˓����^�Y�*ܪ�*����)X��d�h����,Q���k}�����J��kӲK`<f6����E��7��[�r!&�T�0�S��W�9�Kb?��*
�7��2�%6@����S�I>�q�������S��UV���zs����#g�����I]!�FɚOGR���B��i�`�ǥ����;@t�~4�����#�d"we�r	h��;P�Ծ��!���(l�p�6@�QN2����CSyP��CdL4Ny0���}�Q�e-mt�jІ��"k��T`�?��6���K%G���~<��ϚI���h5*4�(�H�X���� 
4��Tݢ�]�:�k8¥�Q0�kD��P�S"u &�$��j�����f&0�_]�d���['&@�;�J�u��U_���4!悑VӅ��'l�i)�@��'��� �^���Z	e�a����YD>�+m��H��q�R�pH�)<"�
�#��{3�t���1%6�i��!�tn�
T�wc��]�� ��Hz�mB�OpI�������u�|�bD��s����2�bU�|m�'V�f/7������� �}kh�
�<�95u?��[�~m�b�4�:��#=�o�]�Ѷ�*�y�&�v1�mo(���(�U*�lt��@18��ۑSN2j��R�AR�ҭ���.�З��B�<��<���SPy"��������`�a�=ihե�����%�>kgI!)0�9�~`�ƺ��Q����d6%���&a�,M��@�q2��,j��GԌ2�|�UŴ6���>�,r?�aT��I�â�X#+c1���$��.(���Lv=YP@Ќ�ĥ᜚E}U��t=:O��g�"��8:�"�jŐ�E��.N�!���C��.7�-߇��d�c����>���"Wi��r!��Ft��X�W�W�^�2�b�H�bPnV�E���X%���p������.s�Hq(Лc6���(Lv��>�_�]�`*z�����HS��� C�>��j��$�����ѵ��v�=�U^i���M�7�����/BB�?��.�nεg	&^4MW
6�v=�'I������X��,����?t�A�|#5�a=��L������'s�lL��p0���B�[�������({����6G�ge� �[bi�+�齓5+����X`\�`e������"^�)#a��EhB��n7~?@���,��xK���Щ�J�A�g��v�>O�
�0������iT���3�-
�hS��$IQ.S��N�:�A�.ӂ?��3�'�"ZR�F��*iS{u���~����ЊX/�<k���DHH�@O1���Ո"�U<B�b��1�+JuG���n׉�gk���`�v$��[J�D��d����ސ��A4*��h�!�Q��Nڇ:��;�F8��w� (��_��W�h�1��� ��߲��*{�U�I�r�}���5E�5{ʮ�f�����J3L��kڥx��2������ћPZ���e^w~I;2��N�5MP���3�Pϋ�T�����߃b'��w���.Xe3��d���G�������y�n��]�jk��YA������Ș������#T)q�;i^�ݼ��M�к����֔^��$`-����s<U��9,�AF��"���7������!EŔ|-���f; 98#Fo�w��I�\�=Q�����.Fk��KF��1i(�Ʌ�����OK�P���4��`���)��K#��n�bZ�\�x$Uݐ��D����á��y,��� ��(��N�?q�
��>��4'D���J���zde�t�C6*�}���
eڼ����?�	��
PF@�#�#�F�Zh�$���ow�+���� R���]?�$Vݺ)����b��h�� ���@iǌŒ���[���n7���s2Nd��rh�eYd���'Z����/]�p�3����uC^�W?�E�2�g�]T}��܂�.��m�o�'mIS\O���F����yg �8�y�4�W:�EW�F�~�X�w��߇��G�ߝ_2K����*��L]��S��ep��a\��U���;�L�}RͭB��(�+�c�ؗ�uyB�iK�#JZ���[n)��G�e
ȏ������[����~���1�J��/���^v�L�s���l
lv�4�
�v�ݦ��ov>b;,E�uМ��퍵���n��IU��U���\��D��]��E�zaP��qʏ��ph~˝<6���K-�}� �Z� �{��;ͼ��+��c���s���:1�GŁ���F���������nF�{Ply�A���T9���
�L��X˨�����d�[:��4��LokM]T����x������p�z�n�4T�{I�Χ<�.2m
AZf���D��g/�W�����娐���_���w���y��G��ۚz�ij�{�sU"I��$�7���Thݸ�B-�9���cW�(�B��~�p�_,��4�g��3����-^|�e!�h��LJ����z^�b][�8�'�������i�
r3������h��#@��)����u�`7���pɦ��j�V>��=4?��.�xy�tAY	��+�zn�v4
\�¶3{�z�����*���\wYS!��{;95_��]	���R��H�;[?�`�e���K��&�*lg�lҹg��ܛR^{�!ҕ�	��0Q��Cg����*OA$�󂀓�rW%L���4e��n(á^�?,����f����dǰZ%+��7�gr�Y�>$���i�C0��2N:K�xQ,?������o.S5!���1���.��鯼��_bF��03A�[w��H�d	V)-�̤�}I�a~<j�C
�v�xF�!�N'�4lZi�w9/NR��ME��!�T`�g Ma�A?�������	<���m���zT�p`-�)��oFfRM
�F]\7�ka�\&��ܕ�Xz=gz/�r��I�ҥ��KG.���܅9#��,X�p�����X��9ɂ��$숱�kfx�%��[LQV	��y �*�y˂�Mc��ԇ����G�+"��y��E��tY�3+ػ��}�D�1�����8�G�<Y�������Y�|�-�4��mu�i��b�3�z�D�C�/%oL'��h=�O"@�'�,�mI���c�~OE�Z^�2��=j{Q(v&�ٹ9�mHU���v���l��-�Ǩ��XN�@��;�x�8:W�1:Q>�Jn�kRR[։���R�/�V���L �N�÷����b�q+�x{��##����n��ClB�#�$p��m%��_�[{�����CW����!�ל� X1V�1�x=��l��^��0rA�b�����%�O�t���y�r�zM�c����b' =o�|?Xp֊�"y�;��>p����-���}VIF�V��٤�"��S���E/���q�|RKG��3�(���"����qd	/If4����W�h�T��~��L���!�j�����S�s�rh�`��D�왮��1��-R�qVNOhu���=�;���V�p�L��\���n�vQ]�Y�O�W8�YP�R�b t{,_��xW~���,�\��FH����)[LZ�` R�,o��uԞa��/�鲮��e�^��nI
?M�p��X&��<D���Q!�V 5����*�����:#�@<h]j��(=���E�����L������8� �#X�$�La�L��o���'��Qr��b�����ď�����\��P0	�.#�f���x}�4��~�sJ�wIhA��h�4`�� �o��b��N�0����Y��)�W4]�K�:`�;�˚��K�0�6Ճ�qZ
{k²��Ĉ��sҨ�k&#�(	����~��y�/�Q��:��p����B;^�:ͬ%n��.���!���}=�$�7�B�3���8[�.]Ø_��Pj����= �Lv�0kaAm5"�^`�0�����O�ǁ�}��ktM��<����B��<ҟ��<J�S��Ʈ+���(/b^���I5,B鴁�8�H�[aXt�-�0�A�>�Q���Ƈ���L�H�~���i�:��������C������N��o�?�{r�t�Czլ�\�/۝3�a���� �8����<�:}9d���"�����$b��ï\o��ی�m y�i%8Z�F@<�M��l�w����{�=C�<��$n��� �܇ '���=��c���J����2y��7L�Vdcз�p��0Y�������(�����R��vỠyu2&���,���p}0��3�W\u*�XB�0
���}�!}���\�ZN���7H�)	�R��`J'a�����ѐ�ci4y~=��]ѩ;N@Λ��J��e`�^�v��C�qΈ�[��_��C��*t^�\�fS[�a*�
�a�gHKxoh[��m�Z�/�7��&��k�>I���B �4OT�u�o>߁w�?P��z�;��;k�a6(g�g$�ks\֒]zt-�?[�m��r1�t�\��,�К� z��!�^0{DB+�!YY:����+�	T��0`�U1��ҁQxJGz�M9E�~R5����e�	�(�LΞ.�a,+�I{y��&�$�«ƛ]�Q@�*�+I���tl�]m���X��c2�����y;��`M����U�&K��50t��G� I~��=rl����wC��%ŕj>yϲ�\�	ASc�G�}+K7ݯ�|�J��8��j�������#��P���PmDdxRG)�"�<T�^��[:Ƕ�4ˌ�{;s5���M��8��^�C1r+cFt�I%� KC��2|�y�?�̿��๫��Y`��DR�8��<����n<��kd���`m	5���02������i�#f@r;g|���rI��a.�c\������r=M��Ŝv��ުsg�c�qZ\?��Ix�.���Я��}���G�#��b��R�0p�h�ұ�|'�'�ʚfp&hϺ��s�^�{��B�o���W��}��B�5�v9����d��k��4%�Fa���)Hg����J��9~�Tx��us�����Q�����U��%����@��L
R��}��U��
��<�O�3�o��lv6�r�>�(�� ���_mT��瑱�إpK��mǥUz��ׅ����f��uKu)ߍHʇ�����L6�`+�U����=f���'tLKkZ˵q�.���'�tx�c4]��t���)�&1܍�6:�pa�B~ᩀ���×?�F�XBK��CH���=�P�yjşfƝ;��m�S���ϕ�#99��'���[���`{$8ssfEm�G��8����{<���f}���s��wW%0�쯬�̔i֓U���h��S�n��6g�hL����K:�P�p-�%���X���]�VHOS���y�>5�z�l
�v=a�)\�2$���ܬw_�����)A��L�nk���H.u�.˰�=��J%�S���x�`���f�'y�<����V�B��u4��ieC�ΐ_��p���.ƣ�%]�̮^!�wR���c�Jԫʭ��7�q�����]D�ϴCX���kj^ ����]@0��h��>�t,5տ��^��*l	s����z�H�8\XV�ް����/�i\��S�fRsE|���˞���w�1^]�}|�����,��`�*���Y�x*��J¤���R����x{J��\喋ow���|M�>�6ƚ�K��'��2v��pᣗ]E���G���Gx6R��}	�����b�ޘ��I���反h�l�4��/�i���7����1�����Ҝ-)��#K
Q��x��n#�LB���~��H{�E3)V
F���7��]1��2mY[=S.�C�~��W�;	@�L�8޸,��=y�D��"�7�K�*[ݒ�*�c��ɮX+���ěP����kG�L^�9���ز��n���J7Шi��p� �_��F�Xr_ϋ��KƧ�d>���{!Ĳ�b%�_��q�D��;2��YY/�N[�}���hnay*E9rp]���|2s+�#�V�'����s��Ry�NY��p%
�V(�J~d�_���(ΑIJ&��ܺ�5�~r�iy^�R��5�
r4�K���ݚ⤻�C�_�ӣA�L�_}�׎kN�C���O5���A�]}0\0��kQ��O��P+��1�|(��T|�|T�-�u�-,�Z�+�L&ȼv$c)��ߕ쏵�p/k'k��#��#�$wUͷ�a��6��p�q̺�9��>�
�%�|m�X��x�_�'`���- l&� E'�g,�~��LGo�o�\�h����O�ɟ�La���'���(��I�zt����`I*}'�T_�3'
㨖ٍ��������o��C�T��xQ��U����'b����'��7���Խ�C<8Gj�+U	�(I eR�wrq���8�:���@�;�$�iS���#�d�%���qw��4��tplX/���w#�P��/>Z���F�e���	�5U��
��I��Jv��%�!J��݈���ba�^G6
�0؂-a#�0?���.�nHHvٹ�����H����Y������jl��k�����Q�����H�fY.=���s��e�@:UQgv(��p��`S��J&�l�Q)[øÜ�ʮ3��� @H[�G_/�k�� M ��Y��,Qpp�<zG��Sn(ψ?�.�!.��v�?�m���Ի�G-��8$���}��h)�
]��*F�z���U��?�*ce����Y�t���7�E?�e��w� t�|�۴Te:�Hy؅��~���E�0���Î�%�ݞ %��G�ٌ�U_�;1e��9r	��U��j
�����}2�,\!�x3�9�D<#|�_�țT��FM)9�i�8��7A�J]°	D�����%�W����	��֓_���(�@T�a~���@[f��E%0Az(�xca}�����h Υ�z�ܩE��0�dQe鄐��a�+Z�`Y��BbAT��֪L�?��'����e�����^(�Uum�}Q"Myl���l�c)�%�� U��M;ƭ��i]��Ṡ�^K����q���	!-�}[�$�ŶA&�?@��>�^���I7����`:�x�[�;u{I��hֵ��D�]�V$�v���vW�5״����L���L�v2i�����m���<��2���E�6u�&�'t!��f|����������}��*�VXW�JQ<���N݀�'�Vd�!�岒����<�R������0Ö���Y��H�U9b�Zh�����b���Ov�G�\,�鵟0���l '���Ū��2U��#?�D(ʠW?p8��S9 㺉x��C���������Z#� ��Bm�[CHm]�O�-#�]�/�B.�ΗW��DQ-�!GGSɻ��p�%�s��@�[32]w����́�q��*������ѱ�t������Q���U�F}v�ر����3{�E�:�a�����N@������z�G&ɶ��t���.}$�ԃ
bix!0,��x�0ľ%M3�ǵ��9Jc��x~�ZX�;��ClܗϨ;����G+$S��p�?�~����0f��İ{r�G������QL�s�������SHГ��� ��E����1�� ��'�,��fY��� �8��"��z�$�=�@����Xr���\�1�jTL�w�,=>�b��1㜇�Sǔu5`�����!���:V��Y��WL[HF�`�������
#�;�M��!&@� y��ϋ�}��o|��&S�OyLt��H\/�e���(�1;W� �.c�8���2z�k�ai�!Lj�kv xJ�j
Q���e#��_BR���Ih��0󝭄��I�#��.s=�o �KN�������@���]�Z�&�C�dǕ�y�\���������pM��~�q��^q��"��@ �%��)��P��K?<����(_W���w�jd�њxV��E��K�'�}���x�	�+j�d��2SL�[u8��oA=Z��$��U ^����'Ԃ��ɇL�Հ�g7K�G�.-��ٗ��[2��c10����27n{���B�]F$;œ��^�T�L[�W�K����G!�,�fe���l)]d�Zjq���ǐ�@n���ϐ���a_�!xh�7�}���� �Z��9nC�z��b�Kr� �7�)�#-�� J�*�E���]bIA]��N������a�(�k�#�+�I$T�X�.�5l�yG_z�>�]�l��Ay�u�͊K���Ҷ�����jR���,��2��)��*TK\aFi���C��:L�<L
�
����-�c:י��W���YU{�+<�K�A�x��H�B���1R"��NN��m���Bg�i�⺲��B��0�&{\����&��>F.M�Rz�Ic�Z�!?hj^.�HpqeV&���[����Te��.��An�wN[�|޶z�/�og��Б�i�TH$,�����h���0k(̵��'N���,��t�gڮkX̌�	��QV�U�-W��P�x�o�!�Q:�<?�9���r�qM���_��\�6�1�?|!���=|x������+p���ڄ)�=�ޡrL��S�KP���Ș���!`�E�}��3%B"�������[b��L�D�Ud���2��ҫFP({K!a"�B��[ʣ�jPa�����ND�@r�[H��j������۠a�bz�~�YY���ߣ����y��9\�F�H�)�"#z���K�#�6��#A���ce]��V�yz~�HͦYy���m.��Jm�^��1��|�쯲����zSa~��].wR��\�tG�|����Y��~�1x��R˳��(���tA���h��{�8UP9R�$v� ka��~Q��i��ސ8����N����m�u(!&E=g�}�1в$̓����L�h�3�G?���+�5!x�R(Ʊ�a���4e�X�t�����3E|&.���9���p�֯��)@�C�}�u!*;2ߩc��yRTT�~�MW�i �ŕ�D����:۶-��qU�M�9� ��<= 4��IV������I����e-�� �z���^[ϡW8�\{���G`��K�Z��]g]̷��Xg���4m��|�����/��x'���R]��J`��8n���D75�΀�(��k�*�_-��I���笿�r�����Mxik|��)�)1��
Ȇa�vVԩy
��6�� ���eGkc�3����cm�T���
5���߉�1�FND�����;�)��^��Ux����.�a��_�}��Ko��8��W=�����~���M���Ɯ��R�C�Ik^٢V���(��Tѵ֧wd�E�v�hk��n=�o��s�s���D��G8����xU�*�0��<�rձ�)�gz���?�f#\��< ��p��4:A�L�;�ґl7��M������B�y�:�=Ն�q��ť1�c�*Åx��t���O��e^��ID�^&���u����dh2�~��E�^�������2�%06�����)��5���r��U8X;�R����K�=�M2�9�`��V�x��ue/�p�p��������U�q��5���x��6XRƧ�����VO��� �8H�o���K�,?���f<�䫵�y��	�Y�R1�k��~���0�|0�[��b����aڄ	��a����ܶbZS���ч�[��q�:��K�	Yg1mB��3ֹ�-h�J_����3�� ����{�����{��4��@�RJ���~��-TN�T�oCC��YK��J$�Z�ݬ����>긔@�m��	�������?�A�37�~eM"x/&�Vɦq�\�R��ͼŴR ����Dh<��ɽ!a5J�_��y#C�����Jw+;C�*�� �x� g��TGqw��Ŏ��N���O|8��D�ICA f������0�b`���@3[hYn��e(1�-�Ɉ����ֿ���S�m5jA�BE������W��XqI�nnR�W]����<O���L����2��p�Ϙ����iF���-p4aA挍#) ��1�<��K$9�8e�-����p�ƍW����o�?ak�0�7)k��%�����Дy�m�Z7]fZQ���i����A>�<,�P�UB�dUV��>��Z�4?�
z�NM��9�}b�ˊ��Rq��aPk�Yz���e�6_H�.]���N�m���4�a}�z��;� ���Q���?�5]K�*W�[�.��C�wx���<|_�%ڪ�NP�T��t42تw��͙�x�~�w��ڵem<���P ���t��D�Ao<����c�S��n&`@1��^��K�i�%,ۗ,$��}�$׿��8j(Ƕ9΄�.�u�V/�F.۪5����:�g6-bFZ�r0��Cv�Ov	h66�ȃO���öujT�o׫��(O��c	�'����>�?��|����E�B� nd�x 9}�/I'ъ��
�%�u��U��}�@dr9��V����^\C��箤�έν�q
0�p�lZ�Ə�Y�-tumZ��[�:{���Ny*���pǇ[��yYyޠ�g���a�\�����R�Y���M�z�)V�o����`�R�}���~8EkK�(D���o�J3ǭ�_x�����fٔ� st�ZF��{xY"$b(�bF����m-h���Qb3�R�����q]5E�	+��P��f�i�Q�X�y�h=gb�BWut���4�Jѐ�ʨ�i�8_��S���������j+&pz� zd�{A��GQ����Zpa�P4���C@��dp֮��x�}���%����&���
�Q����!�/�=�k�UT�g�3���A*Ⱥ7-��D�-1w���â�6@�x;��lE�?)y>�$�:aQ�����V5��֔��d���WXs4w�X����, %��xrX�E7_�xȨl���RTٲ��(�;�l
Փ��?t:�3�<Ə�%5������n��+*����b\]���T�(u�1�Ug��`w.ȱD���N���%R���;~��y~����EO'X�d�?r�IѢ�'���/�(j��E��:�Y��h���&��	�͋����x���f�t�,/�F8H��{��0 �I�U��T�j��]�7Wk�L�W�IP}��9�c_k=X�8�}=3x��(��G�n����sh��v�q��M��<#�V��h�aA��~}�O�s�r�?�]���?�Y�d�Y�f����+������ܑu�8��/*�"��0������K3��6������N}���r%�a�XuK��+�*�*R�:+"�x!�mU$�d�.¯ZΩ��J}ېV[�l�s@u�N ��웨g��T��_�����I�`�n��\������е!jb��"��Ä�7k����VJ��I���[����������U�I��U���������6��2� ��6[�i�d���z�a|U��ֳͱ:�0��}���'����xyH���2L5���6��}Xٸ����3,_=����jj���)�t�{drt�$Q�O=��ɋ<(���_�}W�2^LZ��^�����K�N�R�`�M �		{Aa�`���ǉs�9ut*֒�w4���2�P��E!�� P����������K��8BS�} �Èudҕ}�L�¹{!�.Ps�o1��>��WdR�U��v%�
�y�$������Y��T�;������h�m`�g?��	[v4�;� E"�L%���p����H[�~��T�7)��0+嚍WPM'��"2�l��;�`m$#����Qd/�-Z28j)߇~��!ep!�����Zu3J�[�����,� �����o�즉 ���$)�G*	7 $=���o�m�Ʋ��Q�3�jM�aq����_�&�������M� �19�#)�`}H���O���X��������z�[s*]$�i����R�CK|���P���TV�[�t$T��؃%j+�9A��*�:M;�s��=}��E�W�7�,M_��I������c%���"P�E��}��b��`b����P�4�\��o�:f�l�z�Ŋ	l���@��_���uQ
X�(��Y��>0�����Æb4�=�v�S~�Ұ <�[�㈧�T^��^���6J����@1��9�����X��sjǪ���fj�Q*R������I����<���Sr&*.�;%H<�=�P��_�s4��L���m����knG�q2vK��|��Ig�`}P��)�aJO��n���gL~V��'xY�vI�\����1�-y�J�Ut���/*��VTw(�es-^�ʎou��b���G�������q�_nP@(4�­�/��g#Pk|��o=�9�l�`T��H��BG0ݹ������iAz,�1f�������L�f��af�+~ʞBz2�yٺCaɸ�ɟ%�_���f>6r^�N2zΏ���44�j��ʳ
<�.]��+4���C�a�{��j髰�����j�0?��jB���8ײ���V�6�J�[��?���LҘx����b���#��g��C[]�ZH�#1w�m�*� ��o�n&�7r�gȭl�L4�y7��.;f[b����d���M���;S7t�������
,�5PMRbP����F���?Ʊ@>Z2�mj�)��6���/a>c��7�G�����9�4�:��i	� �R���#+d��͡?z0�2�J�=oP-�\�ACA�W�)a�������>���F��K���#0��#>�="��q�~5��xB���I/��i�� 灟�)��𢪴DƩ|<˔ښ����*�j��r��t�����mYW����x�<dV!�D������.�CG�[%'Q�D���̽��,	��frnڪ�*T���]�|ԡlm����J�1?�A�q�y�Qr�pD�n/�ƊY���|�r�"�z�- �F��Ä��,���Y�Z�Q�l����N��U4ey����f�$9�����Qs��8q���;Y�	�����Ԍ�1w��vܱ��gq��S*��k�m���]�B�#T@$���u��>�?����y�U!�a-$�&A5�t�.�.`�\v����Lx$�o����E;n�Y���z�@�W���3���DZ� �+<k��_'Ld�m�8�l�@�	�>��@�k"9�����R�Ny[3�[���+�!8������E r��!�քn�@-��MHö��朷�J��V�`�&�Gd�-2I7��Sk0�Ӳ�`���<�ɩQnyV���8��?s�,C����k�w>+��[���z	�����Vƺ����5(���̩\ �ܜGYR���]����eT.і�2R(v�`���{m���p��gf`�8A���!�U�WL�g0���:�t�>�6���ʨ�0�)~�����`����w��{K���WзkmQ�^	|�ؗSgc��3Ƴ�22j��K������f�cW��Y��6�3���x�B[hxq�΀%�`��!�IST1 ��S���k%2{��H�P��{���a��������;\v�!\t��{#䴿h���L�N�co1��0��)����z��,����'E��jLt�Q�>��U�/�3D,�6�x΂�v}G��vp]�����2_��&H׋�l�C�y���U�]u]�x���X����
� 9�Bu7�)���4�����'�Ľ�E���\�C;�ݐm��]����짓�1�n��y���(l��Y�}rvȒ�n�z�:���9ut�6�QX�l[��xm���@��nU�ha��L�Q;�!������NPv���_%��hR�bw�[���0�>pR�Wq�l��#y�Ub����ɄKv_��ۀ��i�Q�%�ۃZ��v��[�K��~�bE�9�ݚ��.�?��j�ӟ��"�����튞ZY��>J�����Z����B��c_�b%���`�Fb�:�9Δ�)��q
!r�[��f��q��:컗�#&�7.�L*���;��i0���VHdF�)>��<S����M-p�"5�(���n���>���H '1����o���)\	��Y��1�2�(:�=�5V����M��,�٢-���=q�B������v��q���`ʛ] �a���R��� ->֨t'7r�M���V�JY��A���\<��*E~%C�WЫ��B�����U�̨_:�+_��Z�m�����\��)ѕ&��:�<�A������
R)�>;�)U�T&f��*'�y��`ʢ��oa�/�"��y�y�@�6bq�Ӄ矊��a[���� �ڠ�:���i�D���{d
��5ɘ��p���&Y�	b��H���,ٻ�������y�c�g��4�_�������ie�h2�N�U�Zķ��z$��r@�0�>�?\�	����l�e�F� %�w=A�Y�{��W�9 ���6�sl�����Ǳ�{��p����3�tmH��ZߍsF��FD.�Q�n&��i*�u]��*��5 /?pa������?�.7���;�'�I 7�2A|�4ui���gD��qO_Sq|;�#�4�_1ƥ��G�*��O��~`�gJz�u�#��_�����g���3�Q���pdR��C�\�a�s��~��$��n�0�Q�dJ#}�C	�@�N��k1D�Vo)���9}�J�5��,��C¤�u��w8��q]sX�b��Z8m��Y��7?���bHGM� ��P�����R�1'R��ћ��rhz���p��k��)�8p�����s��6���&rrں����Q?a�Ӣ�F%ןY�p	���h+��Z��%�2�F5sSǮI��`��j�"�b��<�um�y�X����a�N�m���H �T��J�Ng�
!�|bN2xϳ�a*�	�
\�l�>ǳ�C�޹�^�Fʯ�U:d�����SrhT�1�}GP�?�:�["j*ޙz׮��z�4�K��6@��l����"C����k�Zz]��7�3�L'9��6�,�����ה����U��b��ӊ�Ȩ�Xw�z�� �/K��*7"�宽�K���F�4xU��)�n�"S�K��#����&�X�>�+�������b�`�� �������,���lKKݵg%�����E�B2ځ^�8����e
���l`�A#r�5� �����[)aʹTo��E���d���<��	e���G~����6AXc�zk�qe@�߹�e�~�zCȝ��o����qNB����23C�W��t����[[���FGD���Ņ^�/��q��V��������[k�޿�9-@^4��X�[x��8�T����s���~����*w�h��6�&�]�O�bC�<g�ǀK���P�]����qN@ɮ��:�E�2�˳��Jj�+��%eS�>�S��6	!�u�ˀO9��/N�y�<����U�m�F�B�]� e���DƦ$��!ր��G��ʒ6ޒ��b���� ̩xiD�j�[
�`��#B����r���+��n��g�[ �߷ڑ���.w�aTóP��m�@�:[��'j�j���s�
WG��wnt��vT��&���)j/����b� c��c�"�p��	�;H'LQA�ȾZ�հƺh����������܉[���%�&X�c�kQ���0��@�v�j�5�qz	��
���v
����HD?&�MG��72���4�4���c'�$��Z�TJ�߾�{�;1V�Ͷ���f��K:�E�禖漜�M�����E���A&�Ϳ�QV���"��v/m{���i��r�����h��N���!4��F�]��03����{��d�A��F,lLe�]��m֕�N	8�]�" e=\�!�a#�|�.lb�:6U������.%��X^a@�����)��R�j����?	�pq��	P���F�'[��8#.=���3z;|"�c��g�{ΐ /��mM�4Њ�����ّr��"�2xe��z���Ț��S"�J[�Ll,,�EWO�D&U$���R���\G=B�
0
�Fh�&0����'��m]��|+Sa�� �+�]K�	���iWĕU��+�Ә������@�����W�#�1�-�K���IR�՛����RD���}����"!zq�j+� ����Hg�Üc�u���z	D:a?��	�j�A�������yk����I�\M��[�(���#�
�\�}��t�,^�5_��@h�oQ�#��ō��_�Lp�fm3k�bA��L���z�΀�)b��n�4t]�Y«�����6��ʼ~;!L��� V��#�:1+Z`�S� �G}���u�\Y0T����"�B�Ƈ�4�Ӓ!��0 #�-����6�� j���c��F+ن%��1܌qR:z�x�'�~�p%-be-3��H�����!�e/�`�;F�2y�o2����ё^����HiB�@"~�_^:C������܇dq]`�U�V�4��8�E2�����4���W�J���
�r�@P�A��Xh�o��<�?�k��<R#�o�	~�i���(��0�jm_<(��.9�D%4u��3O�|�,!�-a���/�,�9��=�z\okPBg�����+��oux�39+C�VB�Hr芸 ��A��K��S\@���D �Y��19�+>'��CHFS� 9�D_��iC/�K��?j�)8� �w.����QG�������w0��#��Z�@��4����
�� �hM�x�)�p-����g�D8����\��ɵ�壥�`�x�(�K�V��cT���e�G���}Y9ZnCv�dںr�'Z���rlTB�lRa8e�=��i���N[9J�Y��p���L�m F�ȷk�>��g�͛!1ʗ�ަ�'�6��jw�u qo	�|L��X�@~��LV6ǹwc5��5�2'�w��y���8A��%���(�}e=)��!�K�`9d��u�cyЕ
O�/t�רP�����画��U�T��A�Z��$K�3!�3q��M��Սe�'�'�V�:���0)�p�i�i-Z�Ų{!�	1��_$)2h(7�z-�v�߁���{֜i�>��Gm�V!x�hz��:���j��ŧ�e�յesH�'���Q%ai�ao�^�!�~7��ԟĖ�?\���@G��Q�U�1S��ӆ�'ޯ�nk�8��U��eQ���Л�w<�Cq��o|��ؤ(*/`��UW�]�q&�_�D��j2���:�M�c��p����z-��`��t�}�p�$|p������|c��57Vdj�1��j��pA��}�=�4L���-�Ub1��^B�]=_Fv>��ج�qfҗ�G��Y?�i��(���ޔ�GY���N,j@��b`��ɓ�(�&(�I������#C?	���θ���6s�Ieͭ]�W ���v6pL@+��zݼն���O�Ά���X���r'h	��~U�{}��4��k��Q��u�������\}��iQ�yp�P�H���:��?��8��!]Y��r�V��ֈEBU;�E�s^N�7�i[��.�c�E����9Q��h�M~�)���+���W�v���E�����'��f�B��M-x�$��s�/�j�}�5īn�J�b9�g,vc��o�����L�ƀ�Q�$BG�zG1��X�29��5;��Oo?�����/��)eo����܊�N�c��\���Ӣ��"v`9�8t0���Ly�j��F��8/�_G�RC_}�{���13u	��M4�~�OZ�>5�&��*豙���[ ����ִ�����H%�V��ۅ�n�.-� ���#�4)���S@��d8f� {-`�<&�_`��r!��qǫ��n�A>%�49��>b�a�)�q����W���<S�?y�1�Eʟӝ5�nj���Դ�fO˿I�N�+��<S��n��9k�7��P�b,'e�?��{���j�\/ �sd�atRU�Zݮv���W*�=]�����\>�8�0��L����_����� ��>�&t����@�pq�%w�yI��<�d����ܘ�o���<>��C�I~�u�l)3�F����T�N���?�lJ�/������Y���]�`<h}��Ǖ�S�f�֓��V����Â&�c���V.�T�H�>O��m�R�lX7�pQ�ԂP<�S ΩQq9PR��o�%ڸs�y�pZ_T{�_K��o�+t�p ��^#`��F��:��
H9]&��>+/ƕ:-GGH/�%�ޯ���CBt��MTt��Z	̧�p&/,Qrz��WiӒBg@�틁�����[>�woc�I@�:'~+����ESI n���cl`05Pj����Vo�H^6�VF��[ z�`�#ä���=y��l�Ըp�y�5�����).d~�n�u2�Ý1Iz��m�^���"�u,Yk2V�a)����뽯��
�d};!�/���B�|C<h~]Q���L�M:��(\�D��LA��ĦWqzE]P-�A5�Oߕ:��X8`���er�ZUH���෍��#e T>@Av���&�nH�ew����cv������%�jx<0�!�W�����Vz���$������|P�"X(r3�o{�֕ޓ��k�[ZDO��';���pk`6F�5�+�`=��=N6�O��Hn�Na���N��Q�N��q�;��C�C:�����-|8����摍1rݩTZB*�M�p��2��yP��Ze��ВL�Ü���4lO�c�w�N^���0욇89�M��B���d��QX�����Q.�V�^��=�sP��ͽny,R���
#�Y�z03��kcYm�bt5��(P0$�L北���eo�������h�_��l�(v�1�4�}�2q6�O����5o�S��ڐ�|��TZޥ�0tc��Z4^�݈![9E�*���:Z۹2O�V	S���h��I�??10%�Hn=��:������v��D�ĴZ����
*��)� Xt@�sc�N�^S1���⋥�E$��V��d�*��&��f�:��eUL��gߧR�X�o3tT�o���l�����<]w/��}�G~k]��m�k[�GT�v!�K:�>�a����3gH�e�[�[��ǣ���R��W�!���?��zEBU�aTK�)�T���D�J�F? g.wh��Ě�e	�Z��'�;	��F�����s�ĺ�t%�^5��}���
q���怏tx{����ܕnd�(���� S�b�^��5�b��ɉ�d�Wj��b1sa�&z7�S��,hN�0s�~X�R��*���[{&���u�{)��m��x��Y��p��UxC���Hx��i��80����hu!�o�׀��5$Ho���F¼(�qQ��?>ٝ�&��u;���;BS��\�.t����� 4�xM+�(O��h�Ŋ2�IsY��
�A<�?zܜ�)�G��������)mv�j�ᶾ��Q ��ys������w����,۝�A����n�F����2 e�(���ˍ�nv��./���
h��bͱ�S�S�>��?��ṱl�\'�>�i91�0��/�q�m��W@�����X1�sp,��~���)���UD	������2=��Sײu���ol������[z�6�!Ťi+�^\W���9��n��C-��%㯧��գM@!t��
��_rH�bP��B��Q�_�/o���J ��M%��J�q�S������^8��b���E-ZvϽ�	�̓�B9����C���D�s�5�Y��sh�,�б���沖���]��9���"�2f��S�����Y"|�Q9Y��v|�g	��}�p6�B����)�쮋����})t��;��m��S�ԋ\����d��)"�Z��S�}sp�ܖCnً�J�@��fm��c���vqR�.�u���"����co ��m.=h����es���(�8�'�b�,U>���$/��g}J���G�V�������dA6�	_��9ɗ�o�q��s�f�it8G�EȌ���a=��Z�uҒS��[_V~�J5�C�)e�j�:Gl��w�ŷ
.T{�����	���^@$�";3� M�m��E�vZh�v�5�f
���ƸX�h��IaO�n���F�H4~��s�'<0�Z[�vt��c7c�U�7[�-�p��`r��oI;򛰈��U&�/����^�-P$�Pxĩ��ML0G�H����r�2��	���v��XGqS��,j��������O�X�L�Q�=\E@� ��1K��aԒ��H	�^%��TL<>�Ei9.Q��B�N.ü�J�rpA���o�60C�Ř�p�S�S�b��ƽ%��9�+��J2�O!�_�j�)���o��l��� %Fn`��,|:�������ٌT׿�P;�{4�F�� �xK]�j�i�U�E�W�z?>��x��M�S'-I�=�����gq��+��j�8���	/>��35ۚ���XQ�ց��T�N�}��s.��,�^�r@�SA
��h�T���E�����J��O������eM�"B}����ѭ�]���QMq��: ��}A���v~n��Xq� �!FM�@~�n;���+߼۞��o�Tm��&K��/�O�%�J�&�#��p�mx��(�����Z����/�^f��뀡͡�)�U%��Rھn�tx)�]�|dn��J�e�j��>���W��o�&!�M�����4o�0�5:N�����.�R��& ? zX�`8�b�-��ő����KAO��;��=U�=��7���)n��Y�GS����~a�v&.՛}����,�V�(ASChJ =޽�/�u�%�/<٬��[-��&K�Ik��>%�Z:���l�Sd4��=��M��/�Q�+���u�j$�8J	E~�����'��X����-t��/+d۪}XOv_#�R���l0�S �o�rzg�M��lW����I�"�睨P�0O�DYЈrr�����`��N�H��9@�"�R��G��P��B�K�lע)wא,�|)��TA9��5\=PbH�掀Ż �׿��匉:<��j�A뼭�������t?+���{,���B���1p�pP?��0e��_s�΃���������}e���p���Z&ݠ��|�D�~´����S� �-Z��83/|�3���Q�@η]f~�K�������7��Iт�տ9B�i����?���=�ކh3T��ө#S�v�d��5ȋ����]`��;)�c�j���x�{	н�#��m�x�i7��S3a�h@KۇK���rE�b@��F��s�e\��9fݵZ�+W���f��*������I|��=�+ʵ�80W!{�`�Q�-'�:A�k�S�i�nvH1��ޗ����Z$g*4yo�|~QB�����5��O�d�]�gj��Ri{K�{�U��͢�k^��D���/?ts"Dב�]!����3��Za��������m۹����d��N>f!,YsY j}Q;�C�'�ܚ�_PIQ濖��*t�W�ٰ��$���h��
������Ӥ]6�:�)����Y�'�2��(�����b�(L����)#���z�������L�ZIg2!6N.'j#��l��4�!fs��X����Қ.�L-?��q�qf%�-�|���`Ny����]�9
`70s�|�:��Cy�p��N���}E!e�@_9���S��x�P�G�|n�z�����/��a�\	Eحf�O�o��"{p��4���*a�Y^���ŝS���]��c����{DW��N2��2r��;l�9��l���n��ҩ7�dÈ���DR��S1i�M�`�X�u#''-���b�s2��,�kT�_l�G��QD5�u]�5CfH�7�|bM;^Q����~�D�K�ڗ��j�ܒ�P��	�#B%���[ӫ���LC�v�r���+�*��ɀ9�/���o^��x����`|�{)�_8��'B�+a�\>��d�,�O�nKUl�]e\�:��߁��G��pU��d�R�B��Ҷ۷�,��z��+�7��;ۓ`I������=O��f$c�R)%k�b��=(�Ay���V�o������ˋ��J�qs����R��5���
��-z-e}$��m
p͈�����E�\��>v�����@#�3.�7�����Z�U~9*�7�Ɲۛc|�ݼ�_p��m�W�Ҳn�xz�������`��[�Z[vxL>��u������_�jB[���0JM3�`[a?vE�Q4�����łXk��Z�s��a	 <�`�ݤY�q�x7m���n	�|l�pjg�Y��Qj���p�´Nh����vS���`K��d�|�EEy#*��?�v:�1e��9g�%�Wj�4��0���y� ���
"��YƜ���	t�	x����8�u�Wm'h)�['ʉX�����w�Ccʞi:��+2�o�%�	�"�;�$вWF��	�x�6� 6Rr,�%��{��u
L�����vd	e�2�|�6��7~?�����N!~ς&�N�����y��D6�wo����B7�Q�ԳFaFXm���I�s�`W��6W��>K���ϛ�����Պ�D~���N"
��yS���I~T�H�$vK��-��u��N�[��F��r�R�!�k�T�N�C�=��E>ΨS	0�VkH8����iĺ!,@T����kN^&�,�x�a�s���r�q�D	�G�^G��sq�A���E��ҡe�ۃʤ�>k����	Ĺ��#\�E&�٨���x���X�辗�VS?�W�ˈ�L� �5�a��F�,�Y��@{1��=�xٔ�ZS����uQ=����! ��g�	�k���N)�Au���iN�5�훆�ɶ��~v+@a��%<��G	CY�4�5Ӑ�;;����xͨ��])K+�P��f��_��%�F?�_-;N��Mt���<GkZ���[u�/��G#�OZv�m7dhǞh����
sH{�t���_y��If���-2h�>�'8�u9$*S�B@�F���V���9�"?�O�6P�A�5���V�9������Ⱦrh@}���ѫEPdB,�h�spY��pmE�2�:h[o�֎�M\u�������#��Ã��`'
B$]>�MT߰k��I_Q��y�W���L}��C=Ȝ��e���`�����k�Iw<�T7=߂����f��d:=�ٌ�16$��$�' ���s��6vvB:ֺJy1�XmZ;��^�ׯu�wY1\���j0�j�z����x> ߏt���ch��$��R�r@�i���SZ.���i�y��&ȇ�^)7�����a NA��&tt�J�{��R-s�Z4�z��t2]�*����.b�^F�R}����:��sr5]�a����0��79����D�T9WK���90GK!��ZN�2sy�?m.ޢ���݅���r�~'��J ����r׮��,���(^֛����J@|��Up�S���y�k��,��Wm��Z���졻v��F㐄G;�\�GP˄��#�z�4���2o7)��Y����br~���t�vt|�ODX
�x�F|�円'v���/��g�ߕ�w��\������fPe7k򮌆8�c�BW�5>Y�r���f��<D��:�[_
^_��E��~�m��S�����.����g���!И�"��*�*�F�������`^2{s�Ս䢒�RZY�@�J2	��*a�$D��y��˿c���!�
������?#��b�dj�C�|��e�%�P79��p�B�Y�R�cRr�%W��S��~��vI�D[��#@ �n�_'�^���-����u�;���[pE����{h�^�T�c�ӃE����\�%���$3e��օN빛� uѰT�������z� �!d��;eQoq���dJʢt����{�f1�1Q�t)c�|��^/�d�Fɬ��*����<1���Dufgh�i���?�h�U�l�=a���l�,�
G�^ZmO�Y('d�Ý�f5M���������j�HsJ��1Ĉ�t���:�.mV����+S��+��<O
`���E��|��J�x���;�Uk���hjbL��u�Y�r�8͋u���2�E<_R_�d1�AT!�|I�Yё����L�߁��P�Va���s�]g!��Ե�a��c/L������֜h��.��h7���;�>�B����������vQ�J�¬�X�輯��)�!օ�(�Q����^�<4��N���xE�f5���MV�-�*�Zj��5�C2�l;vN)[��'~P"�����|U11K9�[��������� ��gm���/��/+,����wYd��f��C��)6�]u��y@B�[ف��h��h�Ѕ0�A�+��(X�(��:`�f~�yig� �3b��<�1ᚬq�B8z��e�\6��GEE�����G�GE,/�5U��}O����5ְSAoǈ���ʥ3�b���<=V�>\�����{�r���S뻕X�uXM}	!:&�k`&w�د*t� ���? u���;',�/�HSE��.�(��*M30�5r�w]p��#�����Ϭ�)�M�� D�@�OX��T�a�C�=+��yA�	odxg�qa?�Ya�N7S$X=t�YBm?,�Y��f�ay�Vh5��'3/Ҿ���p7�� ���:I�F6��7=��$ڂV��D�H��F����u��Ȯ��\{�D|1��ѥ�=�k��b���|^^p�@��Vv�k�P���9(j�[S��}�i Q�U9�!�TSܥ��ve�Fk�zv�7�h�XZE.�G���xd*[:�5
<p;���f	��]����n�w_A�p=�;e{\���V!cQ@w���/�
R�a��ј[�aka��C�fw7��T�GǗ�X�ˮ�I��n+ٚ�BOa�7)�r���!K;N� ��� �t_I����B��DN̅B����`��s.����YR���@TT�}0q!׋������Ky���`4@��.��K�MP^!R�{2��)�-V�bPg�����2k��'�W�l���j�ۯ5keJ�x7?:9p�s�W��b�׬\W��fX��i8ň�3�c�:��܃`H�m�[�n�	��3�C5��pccP��� KG�9��嬢۶�;w����ꫳzAOH�GG�4*xt��K�PoV���/Ї' ��Ra�n��2h���<5��qi�?u��7�f���%F^��F
�E��0��o�m��,$z�jGC�Gf��ZyR��l��^^���3������!������"'y�6���	^2vz�A��Hq�X����-���()ƴF|�����K�]~�~d��#�=��9�����myqz�]�D�}T�tށ�1X����a�lS6\F�W0������/��'g��@+_e�Xs[��n�(@׺P�EM�D�!A���3V����.%��N�R�/�9	/H�����F v+�㺛:�G��O'�!�5��,c���N�Q׵��'p�(|{�b�bcЈ�|vb�]\mQ}�",�rRn�c&�K2d ^�e�s�6����wB��qNd��6�2Tm�H����z���u��I���~�������u��$�T�ȳ�;�����.<D!&�ɢ�P6�����(ds�R1 U��cW��������Ѕ��	Gi��S�*R`
�\k��}MmxgfB=�3��m:e�c;I7;��hJ|J�$6����֩��r��/�|�Ќ�s3݈�+sF��e1��,tک��"�'�잦��Y��sԫ0g?Lh��2�a?���,@[���J^UA�0�]�,��ښő��t?����`�<����I��9�g�: �����-Rb���f��2h3*�F�_.���TU q�IG�2��v6(.F!u��WBw���U#_���8��sG��,.Q����\ ���#o���h�Z�(���>��벃��]-Yb����xb6J� ��)�ϑ3&VB
W�6�`2؇0�!	_#����"�����mM�)|�A�mv��i���4p@��ބЧ���]{7a��4�!J-������X��z��d�I��픯2{e^[��9��^R�����$[tq�$'5�+��� ���������"}淰�Ug�yB.vYu�q(��Y��j�_�Y�����g�%U�*)�퍦�0�%;�a��3k/an�px��l��0
�ז�����E�#��xB��|&�n��I����ߑ;OhN�	�~�m\t_���o�H�����Z�qu+Vl|$6E$��֖����ܤ�&�؈���P]a�*(i����
Y����&���7�@�!%�:�U���xR�d�7>S�����ӡ+Υ�А&��d�,���z,��B0$9G8��8VV���J�~XY��N*�d�#���o�������wM)Jw�
@.�v'��p�s!��)�/^a�������$��Pv�x�-+����� 0uK���h��q�?#W����A���Z2ڌ��]fE�ۃ}h<%���\��7�C����;���g���2�"3�VR��t�'�a�fe!S��]����PƝi!�;f"��mC�s8��#�h��mF�&��*e� ����)T~k�h����b�-fR%����`%:��(�@�zF���br�,�MJ���%�R��MuO�����'����3�.w�<%
��9�M�K� ���T���j���
+d����u�h�2b]� � S�P��h�/:�JJoH:�����R�Z���J��	k����(��svU庨՝&Ѕ���8jv���풟r ,s�Z� ɦSk�)Y߬)���������d�����B�(l�=a�1�wĭ7��0wZ�Y��2�g�X��ȉn,%��	9| ���Pd�kI+"
���;}�����k������i
}"��Wq%# m1̫�����r����"��-w�N%	��їn�V�묶 �K�ZHF�w@>䌈���E~����[c:6<y�-�6�l<�m��j���\JB��o�(��^���4��7��'�USQ��b'�����ڴ_�U��y����,c_�Z,0�X�{�C6���7�ڳo��%o�w�`2���	�A~0v=N��T~��!w�"f����\2d��xW�`$Ö_�a�8���x4�j6n��`ML*������������ȟ8����V�������4ô G�6|ԉSX����{D�VN̀=�������k6��al�����t�,��"���C�/�`ۧG��{�rGDs�&;����a�{8�ͽj؈�5�	���Wd���Y�o�ޜX�RW_�_ T'�b���D��GGd�>��{T,�����I�.��k�|�H4������O"λ��f6��VFl����V.xj��po37>
�ӭ�̸�dO�����Z_k�r}�O�~UЊ�^�����?�t���-edEQ�H|�sX���ӝ�(|��CHx����ɱ�i��#͙�p/�i|���꺍�"Zj  �y��:��5m'Eﮕjҍ�5j-i<.�<L�[\����H5�'��v�����}������@���i���$�ᮯ�I��T�f��o/�U��A��>�NNY�G�V6�k	�A-ł6�f!�i`b�p`������zIE�ʴ�n`RF�3�5		���� n��SO���F/C�h\�������T�%�󃌊cڥh*��b@����O5��Ȑew��@E��zvE���DT�A�O�v��B*(��ȭ678X���g�j�y޾�2����z�x�D�q�{��Ƕ�i(=B%)�9H��ϔ�A`[]J��K)�!���>��w�Q�=;�t��zWz"L7�"� �Hz�pۄn������^BWg��.����I��E�
�Ff?���7������;�s~1۸����&���lYň	�!<}s��n��,07Gz�8,#|,̭��J�S.ŊN�9Rb��]��/�����z�.���Ki������1�Z�ukdo�7��S��7���݄��3A�k_��G�I���j6��y$0�{�uH�t�FR%*,~f��`u�|�-���M�^�,��?Z�!�����B��h�'��a�e��P�����h��![���V,�pQ��̜��Oe��H�o>�>RB�֍�cٙhܥFD�ǖ!�mۘѸ�w�<��dG+����B���������uΕ��KLE@`��q2���
w�:�����!W�˹+�1���(Sagr�%��[�[�'E�4�O�^��I+2��#[4�ib'?����&����a�� Ē+�KƆ�a���w�i�c�C���=Z�(��Fŷ6b$,�t�F���-�dCP6�H4s?<7�[G
]��crU�R*�0ST'B-���&pW�hVG�=��u�=qo�C	#�2�B�{5	8��_����aH���J�a��V�99$"a#�����Ħc�q}�H���S���FI�$�U��S�e�R*C4�L�X�*,E8N��k�k���٦S<|��+�]X��|����2փfv�>YR�)����OX]��ϗ�rC�0��?w�J��l;.�FY��Bf;B���ʤqV@/kܿ|/U�b]
�Nh�\��)��\���@w�.bH_���L��Y�ï��	��v�-��c�(<����8����Fp������~���5h-��U.DP:A����f֝n�p��/Up���
�C�|ޗ[}����bPM͜���߭(�o�/L��&��];æ�'�[?F{P���}SG�"=,�_xx!bt�~e'�%gZz��jL#�Ht�z�f}��i�L��iEXa��t������L���;M�[j�C�u�F+��zP���l[ATV\^�����H8[BS�0�����PR��a2�=|�=�]�l�(�n���(裁��Lri����1�X"�.�RFiĭ�9+��w��4�?sߖ�λ"MΨHo�Rе1J�\��Ru"�YV4�n�P���~<1��HDK.iK�\=4e�]��I�6�M{Èx��T.�9Ȣ�a ���@��P�y�J�Q����=Yiv�^\�2��Z7��q�>.�{_޲:���\�!nG&�3�l�c�?LF���L|�23���A9Nǻu�ЮUw�^&m]	�R�!`�[*����U]�2�붨*׵��m)�1��0��Qy�9�ޡ�
�G$G,d�QJ,;m<i��E��`\Ϡ���������E���ÙN�JfHɴ5�B�c-|��?�'�B��z�K[v�X1�+�-N�Y[C�%�Mc�/K��.�mc���EPUj9�-�L�t�~(���@�/�?��(�D�4�2�i%~����TDu�
��u�_T�_������;wi�N�- ���*�=�#�G����؛��+h�%��//�<.�����P+"p��_�
<�����|�kLK�J���`
��ܟQ_ ��V�Ѩg��S�O�(�����:u���	5��> Z�w�S��ۜ����_Y)	�Ƣ��Oi��R��=o4c�4�{e?�eI�Y�@�K2J��.�gF]�����RK��н	�}�F*BA��qu�D���#S&w��fa��s�c�y�����Jo�oR�0i<�[��ѯ�?56\4��I�J��V�>��L>�|��n�> UL��Ѫ�}����!g�c�����ah�D��L����q颯)�=�s�N6������I8Щ�Q�����k�u�@J�D�y�����HڼC?��#^jO�V���=���`�%���
s�fR"��=Y��7(�!�|�Sv�/?P��dP�ÏZ[cb�MvuX(]�a7)���������|�SH�I<�2���!��}V� ���mS�%��n�^N͐�x)R��lx,D�8��9�/��߹笻R�?[��3>�T��0��/����I<�+RlI��ko��ϫ[��Pv�&��qm&P�ϣ\��e� �a�ʰ�����-Y����{��c��E���k[Ţ���X7B�cx�7i�!�M���::��cy��:|��uv|X��nĀP������2�DC\�9����얄� � q>1��z�
�
F�u�K��v�b'"e8F	��H����,�����K��'=���M�.x�����X�0���#j��_,1���7�E�����?8q����9�@@�wZͤ��<��:��ؤ��lQ�g�X���Xy�сoJ��Yj=��'I�L����+�O�A2�8�i�j�7��v�}���޺8T�G)Xl��T��wi �d]ZXr�K�?U%t�����6=�@��e1��A?I�B�v`x�A+gb�7\��/�G�FH���;� aQiP~����ja�VZ�t"#�ud�gK��y����-���B��ݢIد�/�������+��T� ��<�h���4
n�[k�A1�h��\+"J2��uc�*���r�x�l)��J�$���oh�Oo�'�0S5�\��Y{h�*���7��a�8$�$ʩW=#��kI���#L6�ݲ�@W����@�b=~+-�-26���S��=�_a�1����R�`�J�zs-�M�]/�����*s.����?�7g������-����+���bjj�����	��x{r��yJ�:H�+��۟;��m�ؓ²�Y'i�Q�F�ƣ��׼�ej�NX�	~'Z�Js��;",Y����W�Ri�AMF�m�nYl������2��RN�?�+�Y>�ϗ�z����*���3Y��<W-N[)�mtN�)�����C�3�,Vd����EsF.�.�����p2�S��[����GU���u���
r��vK2q��N��5H4f��pQ<-֫���dM������d�)���s/�ɨ���z
o�zο�b�Ȧ܃�Jda��>�]\.�[��������)�����fb�B_,�J½����������>f��IX��O�VOW
�rD�e@���>�F����F�VӉu_��0���v"�Vu�le�5�Ӫ��9�[�̴���`$@F+>�?���"A��0��M~
y��^�zsOڡ��ܺv��Bn�4��Y�����W�!�p��a�E҄WM��rFC�.���)j}������W��=֦߰Y�� ���#�5轺����]@u�P;\xd��dK-y������7F����#-������6[\/Ӳh
X2)���RF��T��K�c�7�>�l��%<4٪m���e��:g��C/#�)�[�g��YAzv��Fp�x�S���xg�`B���;�(�I3NPL�9ֆy���
L�X�{(�r ���i�|���=l7|]��`R�"�Y}���<[��Z��	77�l�9��_��$(�
Ђw;N�̌"�g�v6T��,������I�~��K� �68�=cvCW�K���/������w���(�Ab'�P:>�k�xN*��9�4��dj��K��կݣ��@T0�/ z�h������>#XE:6���J]9飘�*��B��@�/I���k
&�P�M�yj޼O
'�f��D��͔?�&u�E��#��p2��WB����?C͵��G��<���Ξ��b;Q*C�X�{ghu8���n��7�.�Jݞ�n�L�DJ�#*�%��噮+�V�no��^���{V���䬄�֠��{�!��.���b������T_8����V�Yl�2���Qe
��ԅ�XJ,*�P.�Dt�y�z���`���M��g�q��`h�A"[�����r{��CV�yֈ,�m�#���d�~�������7� z	�pi~���bE�qN�L��M�f���C��� ������\��7���#SL[����T��h�v�\R��c��10o%0���_ ^�O��i�@����%��AAn����*��u�b26���%OK��u�M��%x-	I�C��`��ʺ�U>�OA�\b�_K���h��ע�b��z<�8���M#�FOj�.��1=�Լ}|k���1x�p�Ap�:��F�r�3�c����cd�+�uF��`�P�U�*K��\H�pi���X�b����A�M���X���e�Ҏ��ߪ>y,��yB��e�H�-ra�7��D�gԕڍ7��=���ɡ��H㵄h$Pޚ�����1k��o�#�?�d[�1���P��<C��.~�&o�
��+Y� �Q�Q$��װI^$�)Buzr~"~	�<�Q ���j��w+$~Y)��>YS���Ȃۣ��,!���`j�˰ƦՑs�%;��3h6��ޥ,(e�?D	�F�ᔷ[���š~��
N^���.��-ް�X��њHxnx1�9ȑ�c�IGa�;W�s&�s;�Hz#���{4�,��UK-w��������K�",�Ƶ::�j�^��X��f�t��j>���ʩ'C+%_B�9��Å�:K��/��	�s �O"<F�=���ff�q�r�0?>\Sf�CVƎ�T��݀ޝ�]��
�e���o���~�5�IS"9kQ9Q�*A�|!�	�E[� �F$��-:r|H���X�E�R�:+:nĠp�l觢ӌ-�S��|J���3K�Y�˒��F/�����O��
��l���bEN��K�k��n��4M����~��fڐ�e������u���S��� ��IdM"�C�x{L�Z.����+`�q��o�ߖ���00�}���y;;*�)ľ��]&�4G@���In�M����أ�n5!�D��;R��H2ª�w�X�St_�� ��S&l����^�U20�ED�ĈI�L���MJ;+���N�1���y��F�������<�6�M��� ��Ef+2���?��P$ĳt5�Ves^���q������A�Ӹ\�qL�7���a=<���ֵ�!n��1�ڛ����)yω�pXf����B� ,�䜊�Au��C��o{��N�2�"TA:�/��V	�}I�v=fCX��ު��5��hK���{�H���扪y�ѵz�)���jNl��~t谼��HLo .�'�Qb�WB�Ӷ�ax����t�:L�\�t�5S��MMq�e��-^�&�t�*#�2����5U��A�t��������|�V�Э(��=�C��6>�pd�f���C{����/7�f@-7�h`#���<$��Kp���e��mt�2z�j���q9=���y_X� y<J8�$�e?'L8>�{<umd}�m�/�����K�"��J��/��%��M�#ݻ)16c��L�Ig��&������khah��Se��cRgiL��c^ؓ5���.��Awl��F����x;��+��b�4h�%���g_]�h�Ļ�1�|W߅�DT�Q� J�:x��b$_�����@�OUD�Ɇb���_�2D����j�{�_�_���
;�:��b�1s�]��o9�?������f
-!��Ƽ9�|�yZ�g��G�A�A�W�$����g#��3�j�M*�����<S�W�a�Ӓ度�t��l��_���F��1`ky�)��u��t5��9��*�࢘G���{���L��r湗f\�ƸDN�$e����6z�&9�K��T)'��I�'4��AR���2�q������qD�����u�1EJ��F��0�&ɕ����Y�7�Q\��_̳�klZ���D�E������MW�d~_opud�aD}x6�\��g94���Q��J{{V̀� ��PL�3�%:-¹�0$A0�4����AS���+�D
��E��+.vȊ���Q��)F��fT�־���<l�tj�J~�
���鑽J$q�HWqv�ࣼ�/�<g�Ttt�X݃��� �~�H��?u�J�q�O��X+hh�n,)H~e.�	X��kbyD�7�T��!k�Ж6x�[$,&Xw]��o�(�Џ]�����w���+�^<�h#��F N�@BU�Z��Mk�E���i�0FV���W9���G�F�r�n��Gyz�p�g�Ia��{ћ����2��Uf�ɪc~,��W�)�=���e�D�_�tO:��ux�A*��z390��
��9�����AJ
���T��hc�s�ß5㳗ᅫ�(�G��'�P@�0��9x��)ύ���i�6�6�."!�2ѡ�N6���h�8���x��2)il�n� J��.���e�pm�$�ln��;�u��pۆ~�!s
����xZ��Ot����'V�&����S��x��*7��G�T��*���r�~r�ɂ�F��J,_�Fu��C���sIU��X��L׹K���&B���F2�i��b�.4�:�OVV"P�0���z�#M-�p)�s]�Sơ�21Ni��2��9+	�T�6T��
�b�m����,^�Ey�S���<b��ҁ���+ȼ�$�J����Ʋs�Y���ɝu���l *��8��s�����m�;uZ�������̶n���[���P�Mn֞�aΞX�h �xD�cA�����x*rp:�-�SF{V���Z��5?E5�òt܎k�+G���� �(5�2t�wI5{�x �����Y�4���}i�|�����G~Bϧ�����l<�z�J� ���_��́���Ͳ&+O@�U�=�̠1�̪�eޭ�W���S��ؖ�� �x�h`誉�,�zwbV��+�D�����-�t���Ӽe� ��~�4���?'߅�~S��׺I�V�!�2h�=�X�bu��MoM�N�M��1�q���[�вsi�l9	��s��$2Ǯ��Ogbs��q�wc��J��$O���2O���f_.W<n�7���N>Y�g��V����|3}���o��y��+M�`�&�Zs�!YR�7f-)����5��;^����+���*�'���XI��R����-�R?�l�D��Ǌ�w�J܅q�=��w��>&q~s� �'��`܎�Q�hK{wa@���:��(L��L�)A�k{)d )E�QIa����ǅ������}�$8G���ȴ�"�G1�C����+��]��lD�ū���bS��lE�v��o��iZ����A��C1��O��t��Oqs[Z�}G�p/`��[���t`��4MhwoK{h0�6�<i���S?��*�� Kٕ޲���R-%u��8= HRvU��&�f����ʑ�~�Cs�Х0S���"O6ʰI$;W��MX@��������RK@.���������f-@`�Ȫ�V<�ؔ'��KE����B,�o��\_��� �u�%�D1=eH����mAY�8_U��%��[�C��w�OWw�j���:ϥ7��9��ػ�aq1�� 65JI�z)�M^~pm�ۻ��6t�^M,��Ib&�7�4��*d�hL, ���<���F/�+}�8;��V����A]=k�ˋ�<�9���Yp��q��%q�J��l��Ai������Ƀ�4�m�q�ܫa�h�0������z�7MPj�k���d\Z�hBL��0l·������On�ha/U3ʰ�`-���Ϯv(o��=�|c��kS}������i�<2z�u�/F�EHNJsr�!>/��^�+����E&�{����,#x�������ݹv=<���$2X.�*A<�q�G���� 0.�"��^�w����2)�����?!���*�ad�{ ?�N��PJ��|2�?�}U
��"}���@b.�1E!+��B��7dͷE>�u��7�f�R$�(ܛ�����B겫N(l��*��-�NV�gqt4z����k�h�φu�P��]9�3b0��<� 4�Q�?|�B!�dM�~�^��tu����h��=��-z��~|g«j� ���6f�Ry��s�3G��)R.a�H��!�\�+)�r��\������DK
��c�A"����d�B�q���[6%���^�,$6Vr*�����J,o	9	|�F����Z�W#cB���6�kJׄ'�Q�����G}q~=g�'֛h��7�V �E��RU��~%�� g<<�����f6�C�Z'��l�*��#{�ԉ��]?'�o�_����}���@�[�G��h�k��<9����	���x�������������xI�-��~���uA�
��t�Q�㹎�,�-��c%� ���䣋���0�iɍN�a����b�H�j��c7�1��/���.^��]����sz�=� ��H����+d���.V!̌��7������VC��M������F�����1hH2���#J��PJ���Q�{ƿ�2��ʞ����$U�̼�������kM���`�.EMM �A�.bx�i�t>Ӏ�-o�?��"am� ��p$wz�E��Yc�T���&�L��i�I��~d�-I�[)%̒{� ��w�����G��M6]i�`��c >��c]�]xZ��A,ύM�2&ކ��W���*^В�2!d�2߁�����l1����d�Ճq���{C�ΊgSw=]/X1����4/9����B�ȏY�̋7b.XG������D���f���a$3*kfڭ"��]t���Hw�q\�
��k{!�r^����9�����1Yn�x�@褈��G�ee >�!��9�:v�p���<�E����2o$��@�ٖ��^X!�!�ksS�
v�A�PWnn7�D{�~�Gy�\q�x��q�˵��E�V��s�W%Z.�C���.����/�,��OfjO��y�DRn�W�Эo�O��f��/��A`����ڱ�1��|�*R�!�YmcP�ھ��t�?�cm�_y�f���D�������v\��A��baF3��Un����5ASUW�;�}胕I���!�Ђ��Ԭ��]��Ť0I�x�B��m���+8�qVk�:Q-�aF���K�[}]�Ǌ5�1�)am4,@�6
pe݌��S�0Ù�u0�E��σ�Ȫ���A;`���[��E7oЃV��0+p}�^(}\�P��ud�9%��l�M����J�#'����g���1�{;.� \dEiHm�t�
��tdE3]�1��ZH�'�6�#j�	�'ڳ����w�s �V�L zð�r��>1�L��PYQ~Ϟ6�5�Wʗ$����D*�����y/`S��>^݌�Y�@��<���Mש ^���:1<�V<믱��6޴�+Ab1�ͯ�<���k��x3!9��[`�>�̧�~5��o�$,/-E[}Lf������uK־�^��^��ޟ���]���/���||����|I6zCoG�k�D7�g"}�w��P��<W�Lw���֎��������F�/4��~z}\�Z��g�D�:��Є�~M��s��B%�3*1E�:n>�,
|�Gc�r\�{E�@�����9���xR��$:���HBSQA/����IՕ6�h���1x�Lb?XSô9�)��ۙZ6��� 9<}8 �.����CI�v���:���o
XWe� �jY�5�rk�Km:J"d���aGL\��j�u�0'�h�ߎs�T��)����zG�Ӑ�����?�Џ��o�~�k)^8�N�w��?�׻�xO�P�6����CT�[g�����{'�=����c���֒m;���;�x�K�&w죈Hb�`�J�7q3�EŖbB���4�ʑ�}�����!'SC$���]�u�ի�JU�ɡ�@{��ld�ד0��?��{l���W?�)˥�5��}�=���/�]jl�8"����k�JL&��I
h��պ$tQ�c�w�׶�^]���5�-6쯚�C��h	�^2B�V
�tzz>���w���^���7Ȼ @�q��s�L|m�®Z�8��a��qW� 5u���Q��m�	pY q.�O{��Ƭ.�(m�IR��j�>gs�W�yT�Uc��n�,�<�Vk�ǟ��@L׊��8eLÂ%�*�����<ϤuO��.�@�'Hҏ6�S�8����D��~>�yyw����ۊla����EF��O?���J�e氫�߃E�m�Chv���� dϸ����CO�ͯ���_�>��H�!	�K:�U�~�h�	"�	�&��~��y36 �!��'�T�1��*2����˱IyeTpH���J�)QÉW�ix�w��j��zg(5Ů�A��1c�;�W�ّ\Cv����/S��+Bn�e���(Ӫ)�mEe1M�i�pQm�ײ䟊��O� �\69�}����D�\��}��b���ٹ���@����y�unF	��^�C��6S>I��zPӶw�O�w��}�P.�O�5�~%�C�C�
�ޭ� ;~k�f3�f�в&�`�?�x�g�H��QN���I�{8�B�������S��s�վQ�Haz��a��k�U����}�g��ee'Qg��z޴
!e���xF��΁����U���&�p�ɷ�@�$�/I;Ƨ����W�����v�	�am���7����4�Y�LTQ��N��U�↴j��Eۧ�~&P��g���7�n��\��	/c��f ��)u���J�SDW��0A��;��3g*�t������#�F����"c	�ϴ$X��<c���������hVPn$|)��A��c��pC��Bzi���y�цUo���d�k����C�"]~v^���csU�-1y��W��?�SF�	�8��d� ��X�t97!���z���}И�'�y0P~�_9@i#;�Y>��.u�m�S�p'WT��Ѩ�Y���0 �bp�����`�@
��*��al\ R���Y��	ZF�4�����(����X���J�f�\���;$�[���m=��x��F�G��� >J3�7$S���U$G��if�G侔5USVD���i�,�t�\�P����o=����h�UԴi0�a��c�h?Y b�>��g����n5���w)>~�zf�m�).�{�u����q�c�N_{"J��E]4g6dZ�s�p�^;�*:�D �L�Eۦ�j��H p
>�����+ rއd��Y8�bX��F�N�3�Z6c�[�y��'7Py۾Q=�m`���$V��-�C���a��q������e����!����}��	�*(@��cZZz��3u�ߖ/-��6���1��6��H-%��c��>I�<�߂��ݕ�a0���7����wsD�ӢQ�t�g�2�0s|�;�B�	���,�̿�\���m(����ǰy�\m��Y<�?�=�lp��7H�@�f��xd�R����@�Y^��^ϙ�ϧ�*^�wK:�dj�%wxB]�5���(�J�-�9)��<?g8�sZ�U���nK���"��MTd9���\�{�/��*��=�X�}3�<Jc��;��>l)ք�3ZP#��bb��&S� �C�:�v�����(9��Q�F8�T��`��~�S:�&������E��A�㺕'٠!�	+ ,F��B�ݽO�H�U���C�/��l�3>�b� �F��)(�E��9Q�)n�2A���j�}x>g7:�ۚ�JW��-.�d#�B�Kj*z���*�rø�m~��byf�	�������1RY�^D�̼�e�d��O(sA.5���(�]_�
���r$�2ʡ�.Pd��ɂ���vk�A�������J�7�O@��U ׇ)�b��F�i�uފ}ҿ������M��:����l86ҏ�]f�k�ة����*L�nGɜT۴"��6>J�Ԭ��H M��q���b|�TsQP����i!0�����m��=sISJp��A�ؗ~�E��Z٨�*U4��zAf��&k����dz�6>��?�@��ʶ'��UI�l��آX��4_��y�M/5�\K��� ���`</��/�!��N�&�b={��vۡ�V�t:��U)yk�l�5R�9�U�)е��x`���:���(Gc51��>Yp*L����ڨ��k0=�����Z�o�R�B���FsK��q�'Ԓ�[�dďI�a�Q��������8���Fu��z��ǃ��w�*�N�+&�j�q�(�H���\��?���\K=����e!�k����j���ڋS��{�2�q���O?��e�a����t��?N?�a�WV�s;�~7j��vw�i9��L�|֓�@�	�3/�j���ן�Uc�<V�O��xk �"M#�0F�eSL���t�_�/����b����7F8�Tb���?^'g��^��U��u�^R\k�8d[��02	n��5;}���=X ��,�c�L���(�`���hl�Y:�G���߷H���d���v�iV(�GM����RNs��h����rK5@���/����!��]���٢x�K�����`�*��hu�8�'Y7���N"�'"@�����(��d�^a	�aZ��C򭣕����q��\c�s��8O��5,���C�j��Z�Y�,�~�tNJ&طg���E0�J�R���L�y��oYnhB%^Wؚ����DW��x���:MHA�9�eA\�����j������B��z�����`�z�{	��P�{y��Y�8i���%�r�A�qB���>ӐC��	�O�z �S�J�ib};���Dh� K/l��"h=���?�^K:2���|Uz/���%�����o��a>�9wo��~��`z�#�L��@Gw�������P�(MK+�Wst�XtD�L<wIJ��}O�0&�ŵG�����)�� ���7;�)�Q��5n ����z��&�˿��R�`F�����7d	e�Q/X]�=��!�	px�,!by�El��WQ�h�
�C|�s�k�fƔ�I �ƒ�Z]{-pM�{��~]�0�	,�!�@:�mX'0�nD�iַK��V�tkʛ{�����e�c�������4d��w(����G�5䏒1w'{�̘x+��hnfis�xF���kh�Riw���\�U�c��fގ�p(�<�i�P�傯Va"��ݣ���\&��E���?5.��y���c��C᠛'�����F��+�9s�'�hWǳQ�-�ު���k�IXP��j�ʶ$�
ݶ�Ẑ]�����B�Z�B��w���E�E�
XnҸ�*�=@�����hT��}����C��pe|L1l����:�!EՁ�դ0z`�B���-(���V�Oel��yݶ�ѽ�X;�*_t��ڧ�6�-0/�l3te:�c�)��9�V��!�h�T���������mH���&q�YQ�#���m�2�[0�A�j�Hdb$r�e
羭ٯo q}���_Z�>M�+ߊ��ғ�&����Ab���P	�!m�z��(K����c��������?�����OW���v$^l!���坯���������C����0�i_)����������	 1�V� M"�
e8F��0�ڋ�sE�~��j>Z,���EE��z4�¡��q��8��n��j����j,J���y�@��2�Hxg�j�n�f������-����U��&I?�����s���N�a�[_�0}ǉ��
�:**�u���-����3�V6�!#�];�#^n�e������< ����}�]Ù���q��ި�z�kh>leB�T0�,_��p�z&��0Ww�n��Ғ��( '�������m�Љ�l`�)���% ��4�-
tKt�3��+�CR�e-`Q`Q�F���b���
���3凤r��^�/h926�a`K�)�:bb]���b��|�j��t���~"�� �+#���04YD������|�����i��Sj\�iaO�jg�y��QtNA�P��"�8�(��¥�ߒ�*_�t�(���:�p,d�z`�za���*���ѳ�(����3��9 Sx�ip-�d.IDS���k�q$��_��}"�ktF�i-s} .��_���ŢI|��1Ñտ����a��LL�d/n-gzV.ʌ�!X��Pm���MK�Ϥ��t�qe� v�o��,��ezn{���D�x�ܝ�t���;1G$�s���d�l� ���Ht��ϺsS� ҟ����{�8*D
Ať�j�����n��Ft�||DvD�	s�M�mH���E�E�.�p�H���/x�~��9Q��)��Ӏ��� ���a�|s]u'D�C$������,b�uj��w�J�	��g���}ȣ����%=\Vg#�n�	yC}�A��($��^�Y�*�KI�k:_� �|r)��vø�7e�4���i��d�E��ICQ)���ӭdFp(��ܢ���
VGxP�͂��o����I�o?��)��ܶݽ�ˢ�x˦�L�L�uƗO�
J�H:��"vԙ����$�υ����Y�����
�����1/ϋ��(���+�`X��\dz#.�p��&��y�
��	�l�����M)Rq��du��&y���Ij�Ϥ/���������Ƃ�G_nX@�+@���p�HW��X����,��O��g�bg!���xײ�p�^{�_�b)�r#z��j<Fg�ɯV�x����XC�s.?�0s��MT��B&�5�Q��!����њP�,�=���1!�JQ�{U�5�Dm�|ú�Afgn��Z�>���G�j�̭�ReA�_j�'n�Q4X!�h���SIa��8D�5�+��9Ҁ�&�sf�*a�oK٘��x�q4�:am F^�%���K�<�!gM����(#!�$&�hS�}�@��2�}Ab�)�!��[3�Ѱ=��WcT����Īe KyO���L�!N�Eq�������	/d��Y�ְ�H��D�,gĀH�W~�JrU��6��H�-��_����+�{��IZu�-��o6�+݂��/����>O ƺs��b>.q�ײx&N�� �C�b�1�K�������Ӻ k���Q�*
�Z�N���td\|>�5-�5��M��mVİ�)�<[�[e��4��@b��
��8z�ny[+��圈Mm�)�c0^����:���U
�,��~��P�J)I�	�E���L�]d��o`�+�e�f=��Xa��W)
3���j�?��z ��ϭ��́\��I��!�@h?(��Fڝ���cR\Q�j�$-�3�ҝ��G��}�H�H���a�[�X�R/�PW��55�:bڥ3�%Z��Pn�2s�@�4��Q&��F[�|�?�,����6)�_�t���,����[��o9a� �d��9h��E�!�W��IY�C��mk8p�r�;X��>:P�'M,�P�0̎YN����Yg9p�|�h���/Փʯ7�/�Dy�,lC��V�	l��Q�hR�-Cn8+�B|nփ	�>��$����,���0>˛=!/p�������:F��W��3�e���b:��Edk�	LI���e܌�C�rF��6q�)��ڛ�D�� ��ojڤ�Qs���`"�n��ų,z5��M�����4ОѮ�eW�I�'�Rkh4�Ț�� �a�΂8ƔњȋNq^ĭ(������U�ղ&���jl���W�˚���W>\���bs�� �7���F�Ǿ0*�v�q�
W�2�ܥw@N9��� �7�3̓	��g-M�)X),-�D8��~s�3.j�s���MU��۽$�*~�a@=^O��{���'���wm=���nD��������eg+O^A������~�YC�u��XV|�`V@?a�Yy��T%l9�����n��׭5��^�(�#�������5�Y�~�і�Y�}@�5h�#��8 8J-q�'83�Mb�A�Lc�r2�Z!���8,���m�j٭��"O|$��X�;�݂,�ϔw��H*�D��|�,VL���>8�����w^���"-U��b��|�෹-�܉Ζ�F��7��'|y�|��,=��,����֣������D�����d79�<��	��O�p�5\�`�;���k����
��������S���� ZC�/!n}J�tK���O� �mɝ�\o*��K+;w�"��v�)��2�E���ݛ&)��^�� }h�3��Rl�1B�w��R�@�_|Dܖ�^*�!�J]��iY���51wd ���P-�+"Bw:�Jo%����Rq_��	f0��o� Z�{�8�\����+�ɫ��eA)IlY팶=��U�m�QqB�5��SKgQ��+Û��,�P£���PC�ӵs����Ѻ�àѹ%˵�R��z<�_��ϓH��;o9��.�B��PF�׉K�b5�u-��H���d��>˂Y?*e�R@o��<��lE���Sߑ��3	�;q.��/lҕ���:!�*�����M=�3Pj�����Z8��KA��ɽ?@wc���g�>��Z� /�l��0DyOq=*P��?՞^��� �b�# �N"�k�A]��dy�������*�������C�c�A�2�b��c\������+b�vb<��b��P�`�<�mG�n|����u�q��[�O�˄~~�·9 ږU���f�S�\caͷS:�������l;᱉r#�3g9������ �i�� d�������Ӹ�̚�N�p�RSδ�@�.���c3�vrL��f|,k2���E�r��g^�e�5ؗ����KOC�\����5��=�S
���|�-�#D+��k�o�0�4k
9_�R�XD� �Ƥc�����d���b!C6���Om��ߊ��ͳ��� C�`����&�d�&5��Wa�_n{���-��P�ݶ�>���]?�W��0�|DW�X�>x!�ܒF�oi]楲��_*���԰�(��p��'�]~�#r���i,����v���T��:�XRM�n �ť������-Z4:'1裝ي�M�Xl���a���j|A^<dy{*�dT����~y��Mk]J�8����;}R]F�/��"�-��Q���[^�8$=�p��E���O#"k�<�xdаM�yQ��,R�Ң�e3˹h�[L��	?���{����,����{L��:��֚!LN��w�W%�" �G���Ss�nP��,��eU|�v��%������x�[>��]wdt������z�*dpPK��<+��(��Jl�+�6_����gZ"� 1�ɕ���2g�l�}�h�}�Y�n�����Q��9��GPp>�=�ԩ��^J,��Đ��"v���-֏��*]��x���	��t޻''i7mB���ې��v��x�����,@�рjۥ��e�X�06�~�b#_�/tmnϣ� �F�Z
#��=���u씿w�#ڙ�WO�k�h:��L��;R�w�{^�>�[�L�1b4-�*ò��ҙ$�u������M�7z��	@H������sr+	<�5N�F����̢�A���z= x*��H$��q�{��5��%�d��8��/�b"x͈��iQ���WSp�-(��ҿ�`�g�]{�eźc4C.L�4�1�������We�#Qn	Hdky�=&���Dqr�1�c8󲻜8�7L_�~w2{D"d�f����%��5���oX���<9/5VA�k�5E��ȩl{��2���`�H���d �&������񠈹)֖�Ӗ�[\�wZrp�r	��wѻ�L[�s��c�+�w�*��l3��i��iV[t�
�V�>�!nJ�a�����߷H!��>��#�>��bKY���L�<�!��j�iS� �H^�q������?�g/��6[�e�ߩw��>�%�Ҳd�T_=�YU�����g)��`��4�r,1G�'53'�#ᚂ���<��]0w����q��̘t���x��X��ϝv�S���v`�v7l��,�mrz��c��9�	&y�T��M�UX�V�{�J�sOS��|��nϸL3�'/�E_Eu�K7���/e��wJ��`j爒���/�&������}���{l(���� ն��C��`E0{,U]%��W�ֲM}O����^d�
I��e�����L0R)?�(���f���*�0&���NX;�BA��j:{�H������	w`��A����s�$�e�<���?�O[a�������iM��?�����V��a3#&����Jp�7.*�
�A�h#99���G��"��N�"�{���'�>ԽH����}�m�[��p@�u	��Ic����s{*g⅝��^}?	�qb]1[ux�U�
�=��c7�U[�[Wz�%`�`˨�6�n�����dY���U���=3E��)anf����F�����a�֮i�]%�Io6��7\f�No^黓}���)�n���+��W1`����{-s��ܳb��S���}��b,�=c�(��޴e�U�f?�������1 ��������zl?�![!����2�C���g�]%�i(�3��/����%nS�:{�gũX��x��]�Nn1'�%�7�9&K��㳣��7����0�{���������^����aʃo~/���ԅ4B�e�UK����5<��4���f7�S8��G�[��r��n����B����OM�)-_F����D:��n1�H)R,\7���b��|���X��GM�d�'��K�L��c�nI��ѱyY}	<�R�h-ź�~>!��!:�x�oQG�d�/0�LF�w�~Y�U\J^0�qE�"�=R��X�]R��m��]��`�>�s�vRj�O�T¿���k��<͛$�Ԗ�=�D�s)|Q7�.^��P�uJ��S�0�x�_iY RɱPRY� 6���B���;�e1�ϡQ���C�7�T�ھ�p��X���s�nȌ�h���)����ӓk]��5X�sN�C�D�,�Ԓj�Ti:O�ʱ���^�N���EA��'�����v��9}~G/1�eI�]v���"�%��j�:q�X��m����$_�>�G��#�����(f9�a������|�iT�)qhf�*��z�Ͳ��{� �f�M��6;e����k��uEx_@'%����S��H�%IS{o���3�bH��}��̠IY=O.'�f�|x�R#�1'f���37ȗ�q�U���\����2u1*�G�4$�̚<M�����vS.����!dȃDdF��������{~�J�;y_P ��>�o�����5)/yn��;t���4�r��@�J	�!�-�r'�\�i���6�,m���I�\�+��Gg��x7}}Sx�i1
vB�\l>�j�luN\�<k�	�OI�����q<b����0���Y����;�D�t�02Gpc=���[@N��5�5���L���HV���B�\��Y�v��<0��
��::`Q]ބN����HX��J*4��~�"әڭ�R�M�bA����Yh�߰g#�y�
���ϗ^�sr��w3�6�p�w|�|����G�Lw�i��Q)�y)�{���O��j9:��J'���u��-@����W��l1I])VjЇN�~uA��Ȃ�8��RM,�<\�O[L
��/[�ƌ�@����G��C�p�Yz��@M^���2l�Q&/��o^3>�w?�"�1�n�z��I��b���˭Iz;�S�Y����߆�p���G������V�a�D��sR\��[��>;ݷ8+@6j����u��S���b$92r	��9U	��4:F(7餤�[���J@#L�����f:X��D�N���n-ĈBLf@�$�a��q��O%��/�2��>Ӈ�w�l�ɹk��i:D��o%\��7LqcmJ�{d���Ҳ�Z�����+�W��zqF�n���=j��%CȚC���H�w��,���.b�[���6[:T�Ι�<>�.������	Q���u!�����Hz�
 �����+_�,/|D��x#a�4�J� �$���q�A��ᔫ������\en�m�
b
P/�ɶ���DS���A��CH�����n���j�u��Ɩ��x|4a3�v*��7�ΊP��.����>G5�2/N4�f��H�!��yFU(XW�#��]C�Ɠ_�i�P�TU�-M��%?��ڱ���v��9yxhV 5����a6�8'=���6�_f9�L"�Y�E��0d�cv�w�TcL+>���,��4z���L'Ya��B�Z�� �z/j(ZwWfn=�"Ft��eVU�vkG��D`܊�N�NJ��1q��n�&h���[<'JH�}2��s"vҴ����zf�a�y�C�h,����ҝ����x!0���^W�{����E�:����+���E��rii�Fg� �}��\��47~*��ҀH�F<l[w�#o|������o�0&�@����X�H��ҡX(6v(����H������t�)�S�Km�����q�@w�9(7_�����j�����UK�cwYa�@���vt(����:5������IR�'?Y@j����ή/��3�/�(�p;N���(�h�5=��,���yV�wZ�@�,�N���~�����g�p�+�P.�l�T��'g,��ѝo�s�l� �����Ը���]��I�z��Wz�޶��<m�l�f���"���;΃q��&C랬V���.���nN!�;�����!���F$y�|��1T@�y[n��[�gNJߐ��pD�`c��!�풲gk�qMF������se�u) ��:����Ӹ���0��В�fV76���ȨͼVu�ҹY�j5I�Ro�p��~�Fc{I'�wj�E�����[�ӨM`��==�[�ob����뙻����>E���?ӟ�@Z �A���������Q'Ĝ��N_7���MMVօg��j�^?Vs�����5z�M��\ݺ�jd�_�?&?}��cWD�;��Z_<�̜�;��L�/�yڍ �[�7/
�����������,2�h+����r>}2r�p|�t�rL��q������S�S�]3�(�͜���bÅRg4��`�`�{��&_7K���Z���)Z�f�ۄ��w����A<��1�K�ED��an�x���Bk�\I��\��?�с�L2�%׾N���t�SB8��Pv-|u�C׻jH���Z�x�#Ĺ`��t%�3�gr4*ʜuL�΅U��1��6E�	��HB����Lzi�Q4���K���"#Xw�υ6��G�(��W��N]�}����%�@�HAY�9��p�D�NH���D�S8]���Ve�BKjM���&=�L�m�7�L�����ot�����|�TxE�%
��%�H�ºD 5�r����q"�֓���'�����ReM ��@ρ�V?ya��~#��C��Y �^N)�7�,�|j�.`��&��f � �7�f5CA�"W�^R�<��e�2�B�j�9~s�ݨ��_K�kdê�
�^��gT�Z�F;R���
� �Iƞ &]G�D��҂�e:(� �Z;`�w�m����C=md��@�:�Le��;p��n�QcȠ$k�P��$�y�:���g�S���1�F2�����2����8y����t#`���I|� ��-�펗L^۱b�sиu
�F�;?��g����اW���	ܹ�T�<�qQ@�g�j+�m�(���Lz��C?(�'�yx�Zi47��_��Ռ�Oج}Q��BN�ƨg,:Ԭc ���Y�"(r����'�Z�ٹ"���Iȡ�!�7��.A��w�ln���n8"�{��?�=�� z�������E�酩dNNLBk��PO�Nk�t�[+�AL��e��F6�/�����n~LJ��!�j��d�Kx'��b��z+T���}]�r39�n&5^AmW,#�y:n/��ϥ&���c	���)��
Km�U�\ŗ�����Mр�$xå2��'a L6�j��n���1H9��7x�B��� ����[e�4>�{t(���`����Rɽ^ͧDUh;�8ˊ�+Ť�ub,��L��ԢԾ#�a:(�WK�T�\Z^u���Y�Vk;�1p}�x
A��B�CXk�0ґ�\����lk����B@e"��H ���q��s�?{��Y�̨=��ں%�b�?�������=���aA�n`��E��~�n"#N��Ϛ�Ч��N�&{�K����\AP𠊔����/���P;H$�)b���z�ը3�k�ݥ����������	�-��>��턹�[����"��R#~s�hi�N�Gҕ�.�D�[,9�GY�S����e���ѭ`)*_�:{�{A�;k��Nz�a�`�%�3+���#���S4�S�n����&w���jf�j	ZBN~KL�#���])�B;���.ƽ�"%6{j6�V)��Z�˧�V%2\[�p`)�D�%�cq����)���$\9{f¬�6TИ�F3<^p�;�\�zs�=kܿpɈ�&v��V\�{��G��:%�&��n��O��	n�!�K����g+o�!��z��oR�^����N��5M���*�%q�l�p��R&������ɑ� �W�|A?�ߞV|�>C6]!]����E��l4]�g�i��+��q�,��׿��ei&T�b�eD��_`����僣8������G(O}�(����������)�O��5����|�	�h��%��h�Y��"%?����0�����;�eL�N���\g�K�ItU�}MO����}��؎Ke9I"M��y�;���|�"�5�%g��4����2F{R����ր,iSU�U�)eKw�g�
�q�����4��bO�����T��pHw��=��9<<܃�� h����9�#~x��w��,���&M�.�,�D��h��O��ݽ����_lq�/1�?\����o�t4l(�(���Ӻ���;�1GF׋��F�m#[?
-�(F�&*!]���@��S�H��G��1��oc7 ���2/1�̛C[���0]%X���`����� ���+��s��a$��0`[��a:�`��g���I��$��0;���G;!w��N�MV��;�,�	@Ilf4�UV�����'��R22�4�9��� �}o���K�5�� z�w/de�:Q��rßR�=�p6?�ܭ�7�#CM�����]r El�1e&��&8���0+;��o�V6k��EG 1b�B0�-�#��<#5�y��@q�	��$o�oD��e
ѱ>�C���mj�]���},����ׯrz+k�iј/XiF��H*�r����<��E�}Y))&��Ǎ�//I�Ld��w"2A:�F18���{��q�	����gɴW�s"�����z{z@���i�\� DU���������e�`������n�F�@�M�L�����.������u;0{�	��Q���"8w#[�A �y���m��~ޒUѼ
�zA����A��n泰�$T}�_��<�v��FK�/�Ny��xr��ܰ���|��A6�����I�K�#B/q���*����!N����A�!�Z���aCc�[�D�� p{�3g$�D�ctd��M�
�$��&��~XT��<�H����vƚ�V�e��A��q4�s����
x=����4$��P@A�S=`XX׀���Hb
����D;������dXo󄆀Nn1eX٬�N�J��HO��U��g������X����]��r��*���ؗ�1/$��|R$�����$0+����@�k���n��S��8���Y]o��[r���s������4D�,�u����S�wn��4���s��Α�!	kT��a^\���S�c�"ī���D�i��Y�	5�p�!ت��{���5�$P�~���n<u�N��_K������H��*�[��ð��һ[,�!7���3+�9v=�����H�Y��=X���p+��
p��y\�W,�x%7�(�t}@R��}7vk�]@rf��c��UͺX-�>_�v॑���v:_A��=�!�2(E�8(9���3��oߵ*���*|K�mt����v<�J�j	�M1Yϔ1��$��Ȥ�=K�~��<f�؃`5Y#���E	�����[��c��7˗̗�;}u���f::���
��F᫊��.D-u��t�;%�j�an��Q��<�FYPuZ�Y|�	�4F����[�!�Z��}"�x��E����y��Vid������5��	�"�"�Xك*d��E}�f�����-�����	����i�b��I N?���80@����:��J�����V�&<�f��̰��?�#���$���j�쿎�?�_��w����	̗�o�d�
�D?"��+cW����L�u{ta�Zvrw,R��vR#y���!V'���1z��rw^�֦�AG���[P�[p{@֌D�{���K��u[K��T���D�q�S���<z�w��I.����Z�b�աhx�/�_����{yJKW\b�1� .w��DU���dP�v�	���iX�u-����e�c���	;�
'��
wY���Y�eJlt�lG�K�G"���Q�����$�D�j���Al�M�6}ii��1=��E_R�Ѹ�vj�|�<`���L@�%���s���f��70�]�A�>��eo�R"��Os�J��a������i7��0[ֱ�o���H�V^�
�"�������F�FZ��&p���`e��H�	���K4M��%�����ɦB)�)�A̔��"<$ء��!w�ڃ�
���0-N�|y�1�i_�飇IKCi�a��8��$����J�[�I��{�<xvܞ���A!E�ag��eI�زc�<�&<F%mJ�o��Z?����iƼn�S���x���_���I׆��Z%cc�V�5Y<�c+��$m��ax!��8�'�¬+�٩^q�b��X�e�D�ie\7w��K�vG�8�s�; /
�n�Z�
���� �'�!�nʎ���ct��fE����u��'�R�\�� ��K4ڵ�Y�f��Y�[*��w8��C�!��,��N/c�����i�B�J�N�e��~�,
��^/4�P_مP]� S�5-�_��$Nb�qdw��c��a�f(���:l�~��	v���Ru���uP�h��v��(5��O%g�.�$8�X�C_�l��9�mVw&��܊�B��Z�HLM����V�@��&�3�)�nV�����VX,�Wh���)����*q)UƸ�$PH!�R��i��G�A��)o3e�e��f���3��U8��Ⱦ�3:�ᗍj{@���]U���p�b��r��!E?w� ����u�'����m]N�*6(逤�8P7k�ߎ㛶<�I�W���:,Nk�ۉ/	�����9���w��0Bv)���F_����Nn�wMIHo��1����Mzs8P�~�)'�9������j�߳ԭ��tT�R������ʦa��G�O���)b�'�K�ߋՙQK��j���$��6A�����J�P�H5�����J�G�h����\��
g͆��ȳa�e��yJ��+��:(�y�����Y�4,2�.�ACJ��",�x�߂��.�Mu�_�kx�����Ocq���,r(VEy_|\� ��b/�c�P'��l2E�%�� ydR1}_��/�e/з�H]zȍ����t���]�农.���aq���ry�9�5O�f�R��0]�Kbo�)��a�K�Y�ٸM��H�@㉝h7X�j��_γ�b0g��OR����P1j
Q��e�w�Mz�'�t�kǀ}P�ė>������U�׺��1�X���d���A,�1f�ʼ�����|yXH��u��*��:�'��O�ˌ۱�� �	�!e�3�������a|�럯Xť�'p��%N�C<%0"�Τ�J�(�a�	-��{�:6R���	�O��
U�G�Bs�c�趛Ͱ�w��f��B�5!,:����?�k��M�Z~�� }����ri�Z�ء�~aXl`�cl�G�T��F��z[_�վ7|�.��M�NI^�jf�V��[�R��L��|e-l^`�n?��a���To����?#�O�n�1�+<��2��SL&f`���bD���zW$���v4�g�-�1�G��%{o3��+�u|}B�%�g>�e'��tV��쳉Z!��S?{�Hx�L�ӽa�[�u�ψh�m�z@��������w��L)���Na��x:�ͳ�ষ>u�SR`w.����ӣ���[|��D�-�Y�ч[��++*�q��p�'�_xX2�#w�>BU�)���Ű��N�=�Hy��9x��D`��+��'����{��'������Ϯ-�����B%=]̐��f��jr��4�H��1P�bb��~Z��U���0��F܏��w���?<��[7L�0��3,:.�Hٱ�DN�r�ZA����/7�^/���P��+ll/��JO�À?J�)C7!	*�o1����.U�BJ�5";���E�Pm�z��~Ɇ�����
���BN����U ��Y�-Ѽ/�L �1�<��y9 ��|��V��]��	Lv�Y�+��L���h�`� �>jD.��#?�jO����,��Jn�|G?�i���tfHd=��_���ϜMR	�����h��k���.# �P'��v�O�mԞ�����t�������'>��kxo[�wR�)��K�+�t-�>�]�����4V%�	�ke�jg�W."ɻ�X���T*���/����n����d�44/�ш�;K%$�^�����a������D�����LQ�����DŊ���V�ն��l;��Ee|Ng��ۘ!�P����w����45+&}����Q�]u��b4O�J�������Q�:r��� ?�ͭ�r%V����w��v�duKΐ�T:����H��Q�ko�����D6��C�.��c�3OC�#p�'��x�c��
�k3r�#.ӂW{z`�Z���f�}�<��y�2�\D?�}����"u����t�͑�JU�d��ݬ[Eӷz'�J�-?2�����c¹
��}�{EV�Tә�D���W�Ü$�9
�=2��u�K�<�7�_�B��U9<�q6G	e���"�9�З�����x�����&�>�wN����[nKH�(%KW/_f�M\5Fc2�^&�7��*��zo������H���-@Zf�x?�t��fm�v�m�S��?8V	5�����B�od#�hZ���0S�}BN�ƅ���t=*9dH�9F����7zF�6�5��;����Y�h�1'�?��Mͧ��`��s�Q㰎��Z9��������jnPbc��M�vsk�['~��p˃����U?R�`�/�~�AGl�����PeC^��Fʅ��G`ޯy_�(�8Rא� ��B��5}d�Q �-$�V���\��p�@� ̂4+��#��D
ԏO�1^���YCu\�N�^P��1j@lU�v T�|�����j!��	$���_����'3hY�ԉ�q�^�?�I��o�Қ�S�O1W��[��V�~�v�����O�!KZ�p.�}�I�����v�U���v��*�σ���dD���f�o�g��|�wK˴$%�	Q��;�#��>o���{0��uW
+�JC��0�'�Gȗ.�g�d�*�,���6^
�� ���0�����^�[����\��� Z�v�O��� �(�Yyr�'�7-(�%3�sR���SX�2��!��0(�M�	>��'�����Z�f8��"��t@��_�K���&�+�Q����/��gN�����BH�<�xW��S[�D�����a`�LR8�'
�H��]���2թg�F���&�w�a������sj�j��6�/Sp���ltq7�A��v@�9��I�Z2Dm�^���}6��)�����Ĭ1����(���[�8$���(9�6�`Za��7��"RD�����Ѱ��<

�2a��H
�2���L���\��U�a���p,��!�����P�	���D���F*��{���S�P𤢥�L'x��y��Q�8ę��W�i	��-���tq��]�BB<�sq*$��%F�'��-ez��N�w|r�f���������L��{����#�x�� Bi��{�F}�?q��2�����0ps����,�3\`�lo��1�_�H�R�pBOgU":8�2H.&�aL��	,G�QO��L��t�Dk��Wߔ]��D*�m���8����Mn)�I�ȋ�_h}�1Aq�(hA�ZI��p�P�\u2��P��i�S$���ۓ+�g��_q@(�b&dh���m���_`��/dǲ���-���R�J��z���+���?����w���7���	(vN{Cܲ����Fw�i�643�p�{�.מ��!������mU׎��s���؝S�w�Ø^-�(�@^��8�Z��Mx:���čE H�JL�O4��1�oq�9yW�%�cs�iX�-=S�_�z���e�Y9ά�l�9�L���ϯTˮ���K��&�4j���{�g���/�
�|~���	lGS}O�t��t쯐�i`}!��b�49����U{"2f��|�h�!`F�����,|�ai8�eh�tzFg�?���S{�S4���V3�"5��iJ_;�) [�ʹ*i]C*܆�y(�,r �+�/��ӛ�７WH�nEN*����,��j�X�̦���VG��F�X�$A�tco>K|(R�9\�1 ]d�f��(/�.�
�{f����*�O[U����mBX���v�y�gd,W�|�ѥ�sk���?c�jU~� ��2s���nl=�Z@"��c����f�ou�� ��ș�U��A���։>��,~2緙n��Myk���
��B*}��yl����<�v��Ւ`�l��_��Ɏ���B���8W������pב�P��.��hW�����>%ݥ�Y�e۝�2�d�����q4տ���|*{,�C��j�E1�g���[� +��6A��Bq�[>µ�|^�`%�cH]�:�ր�����>�e�jb`e^�÷+9mG�	=�ws���l�����9�>�n�ZJp1�}�RiP�9.*R.)�F���E.<(�bt�:$I}�{��	ȋh��R�����p�k�3���͊�b���A���i)���V)!?��t��m�Ü �<�eW��Y��6��H+�B�����_�#^&�NE/�����ǜ�R�AΐIܦW�T��}�B�$�P�0��&.��
���I���Nv恵�=������N����E7����$��Ȳm��q��	Tm�rhȮ�5�*������l��������}�n�I�-k r��u?�9e �`(��z�(�=����iР���ɌE�{p�$��d�'�
AE�1X➇{���9ҹ���5�/�Bؚ�%�1K()vJ觾M�4d9+~QV���q����T�EH��q>& 5�=�x��^�.�k�a��9�o�ŶR���1�L�SN[29yR�o�t�8�+)��l�-��!��%����F�S߾��eA%�*����g%����Xy$\�{�ޮ7@R�kX#�愨(��'��5�����Y-8���r����C������ҁ��&Gw��w��K�Z|#h��\�Jw�V]�@q��*�la�횀��F���N��_�]f�
.J�?�i�k���>0�`�ws���y*o�X��^�����:���E	��H�?"�qz��]�N�$������V�Y]��M����K��\�b���>��!8��9�i�xsL �a<s�K���R���ָz� �� �z-���" 8���O`������)h!���?�).�<��ME���Ͽ*t�u�8�t	D� ���E��bD��X5�r��Fo9%�n�<�9c~�4>(����ox�D|g�r�h-߹oys.i��싴Ϗ`��v�?Y�ݑTƬ�5%p?�8G�)�(��vtzT$dR,��@C ӈ6���Unr�NN�>�+�|����Q�p ]�ǘ~�����*N$�5\nG�գ֬����Z��[H��a�ך��N�f�����=Y^m=��a������6���#ڰ�r�~oudrn:���֌6�nUFlj�F5]�l�^�]%�Q��Ë�Nc�����[Y��R;�M�6�vD��� �kq�jh`n
��1�sJa�N.�z��]�ޡ_���R,O�V��|� 9�FSEuB�)0��T���q�������!�}�Ȳ�Q��G�Ό��.�=�+O$2���8��92&R����?H���2��4���P	z�b��n=НjP�:�l`�wxMA��M,�B����}�ׇ���.S\��<:�?��r�wޱ��6|F��|50<W��;:�gި�+ 3����Ot�&��g�Ax��p��͍AK��y���CG��U�O�i}��1X��ۊa�<�,��,pk��;�Z����c������v3W��OѣFu�ؿ�Zۯ�R��2�:�,=���	%�R�U����9���-��i���<�q���Lk$-g e#�z�u��k$a���sqg�Rx����O��R>3�oѾ�O�� ��
�3�����bz{�7����2G?<o9`���rs�X�QE��Nf��!l���[�J>�WKT�OH��pj�l�
l�_}3�V����O���zd̊áɌ�-��`�O��H�l���JN���,���IpA��&�֪�O�K3 ��Wyo^&��F�t�t��ω��eEN-��f�+J� ='Xсү�%՘N�
�(D��������0�j����vq٤�g�4�Z��
�9�B3.� ��q�ɻӯ��e�� 	�����%[�4��<:���:�Y�O��0(���(�ɉY3j8z*����pe��}I��BΡP2��M��2�;;t�C��9����'�Cso��,O�ճnU��g��ZIT����"]���&��2s��5,��6�m�e�Z.H;�m�<k�r1'GY: 계�ŝ��z]t���?gu���o,u��z���}�!G�/�.�_:ɂ&zm��-S&g4MTIq��n��6.]�y"�dXo�
��MvxY�B���f]ϷZ��7+���@$B�/y?�y�.�f@�t �f�-D��c'��#ܡQ'Z��{�.>+�w�A����(YNN��Й����p{j�5����[�ēȇ�ē8;I��l1�:󐪚�'L��n'�i�tG�ۀ��S֛�;��]f@PU����GTR�-�'?��k�
U�����f�|��|�p�ZD�eF���?����h���U����>�NK� �qЅ��;kr*>@Xb��iq|�J�E��E�_�c�n��SЙ=�����Ϝ�Rt���,/�Q�I�h���&��I��<3	��X>WY�$<X���ٖʘ�!������{.MAL����2dzܽ���6�6�˾���TE&��q�@j�g���[������1��]������6�y��e�:s �Ż%�Op|�����[j��ރH����(iS�ǈ�0)��P����C�z=����l��;hP�yUijx�³�����`��ɢ�8�3Q
��k��2)U�;P����� |��*�m&jL�rq��H>�"�!j�y�<������C�A������v }Ta�O�[�A�Xۙ�Lg��H�+L`�o]��}� �����#eD~�]�i�*�Η�!��z��,�����:E8!.��'L�D�����hO2�ٵ�=I�	����7���S��4@I��Hr�����L�oA���mV������,���B�˅=L
��R��\PK�B�P�xޠ4O�E'�x��	g��t��L��,��3�+Nytuff/w{�t-�J�NfP|���6��SF����M+�͕��,R��_���W��*�̹�������e�&} �"K��.Y���=�8��K�6��ٿ�f�5��]Z)&zTc��~���k����;��d"7��I�
0��-�`>Vt?�������9�tA�C��	,,����5���
j�4Y�g7j�vG�d��O��9í8꺅��s�����!��0^�vb�y�j!��w�kp��1��C���=P��/& �f��.a�^��K��M�.; +'8���Ld���^�u���m��Ld:Sh�4MN���pq��A%��n��w��[���3߸�P�A����+Z�`y�B��:g^��h��&J�eá��U^y�j��c��I3g��Q��m�"��NV<����	Nx�}�uO|��>HP3E�cّ��4�@���n�zkљ�ۋ�85$h������R��=��+2ǂ���h7RŪ�! ����9�܌�Ue_e�s�7~Q���O*î��PI�\�NA�"V���-I��m.�P�7��W�=����5�tB���͸�S��%49ë^�_���/+����J�?l!5?�\�-�X��y�}Bo�0��wMV���m��P#���v�����d��A6�
�ȎDV�Xj+��Ӱ��H����2+V��5e�d`���E^r3UgE��h����$��a
A�Nz�.'�BE�g�o���Ca�(9�y���#�1 b�^f�%G\�vC�uq#��A`���m}c�!V1���/H�H!w/�@�K�����ݲ|������'b�2�U�w�,(1_o��&]�Uo��%�@mڌ]@�ƹ.�~�Ԯ����)�<����ұ���?BQeB�����]ؤ2��u�����ڻ��C`�Ι������,+��o"O�&WA�E*����`��X��<OO~0�#��@���{!���5����1�C�`n�O'{������ ��T���E{�_B��,Q\H�{���x��P�t��smf��2�T��qѠӕ@z�Q���	Idޛ6��)����{\������� l��:\J0�<7V�覈J�W���w��.{�y�n���n��*�2���$��}�$��"�`�&����r��8�|n|�A(p��T�N�,�g�� �޳ؤU �l�Y��|"�;m�kP.���>{�;����u?�s\y��2����e�ԉ �m�?��+�{i�
	b#�jq}�x�����?�>`��[HD�l]Y��$h�v�b)�y�JY�b��Ps	!Z���� Խ��hT8D}��Ɛ�2�����w��t�t��@�u@��+�E�+SM܅�m�q��
]`�y�Bc�n��.�|J/��lB�+4�w�᠂p:e�+���iE�J��.�})G2ET�_#�6�;��c�6������E"�׆����mP���4�YC\S����ˊ�W4�0��ڐƚh�K��k+���gT �����fQ�D��ah�V��@H�A�i*�[bPF�8a�&#E$Z�l���� �)P��i����8��?���[mPo�X���W�l��ٺ�"���M)٨���G+��T���v&9SU������,焩k5��;��~�R
h����.��6l��
���U��7%=!5|+���L̿�`�����m\Q]x�'c������އ.-+L�귭�y�7��v���e���#�\�o�"wD$�a^�)�-!�t�Crn��Җ�x*�G:�i.
��HϻV-S�[fOg]�����t�?�!�Lo|=�V#�h�[�qHm3>�D�bG���C^]�Ŝ"�5IAGơF�G
Z�xeJ��� �����ϝ�MUl��16��H>�����Z���1�ʁ��k@Y �Wӌ�R�n���?e!mNhS��{@k�GQ4�ç�&�3�&P���hs��A/]��k0��D�Z_�+p�L�^�.s�o�f.�Wx\�f�}Z+8�Q/z�_2v��/K���~(�'�d�K\T�jR(�����*u��tl'n��~l�8���<���v�p}�\�wN�M,���!V^����fVwؙ7�����L�{�#sXk�2��1�Z���e�(L<�B� 4��Bj�#ū",�t�pt`�wk̟��I���yz|�϶
Ĝ��Ť@���/��s�Q(�V�\�z�~��6d�"��^;�X��=��AK#�ě����D( 7��vS�x���"�GX��A1A�V�tI �@ݏ�^�ꖲ�!wO��I�_VN=,�O,1k�뤨8���PE�w/8�~H,9�7�$Rw�Ȕ.i8�B��d�CP���4t��T?�T�+�����qMm�w�,�&bS�^�7��U�l�!-s���m!�H.ՠ.����_+;�IY(j��,���?@�h)���*�!Q���@[1��QTǼ`ʳ�#��Bw���$'77Jb\�Wꉄ�b�ZJ�$�q�% =��[�C���#iV^(wm��Mڗ�z�W�=�a�0]�])G�O5c�*��X�r̰T����K�A���,�
��?�f�W�P�\o��[�1�� MuQ%�Ho�/��p۪0��ZHMJ�Z�
�V���X��F7�����OF:�E�M:#_{
�9��Z&�'I�iv�ּ��&����m=�Q���mOX�4v�Cd5�t�}�Q���=c�?G\>N���9&������7_if��p��.�TI&Q� �F�Z?� �03]u�b�A��,Xl�Ū���f��H�Gp�|�B1�"� /V|��@�p78����}�䯥]��%W�K:���x�@ n+���EA�iV ��89߃�
������F��'�B���a�hw4ņwlFX34����>�4������� �0��9��]:d�{�J����&T���W
��ܖ7��q��l���~��+�6�}MI�����xVr��վ�c���'z}y�˒=j���<V,ȁ���sn�\ټ9(���<����r�y����TOf6O��]z���`n�p�"����u�Wa�0-+_f�0����v���]1WK�Ք?��sא#	��ӏ�0��B���B��M'�N&��S>T��>���R��#._�ծ'�����ߕ6}A���
�FmˊF\�(!���è��Ň!	@���s�+�\�m�9��E34~_�bՈe?Y�ܤ�k��J�LiC�^�U����4�}�C7��D��pm��i�<Q�G~��nw^��.>��#*G2 5W����w����@���.��&c@�)�_�y�}ҵ z�a�'	�,VLW��<�sP=�~�����4'��)�
�q����iuez���I�k�sk�|*��r��HE��_`P�݀�!�E�Ge Y�+�p��k6e6�<%�����It�IjD��ΖӘ���
=2^�IM|��Q����l�~�1�:�	�Q��L�㈔*ȋ�t�!������=?��癁�j;?Q?�X��_)@8i�;���R��\2O�i4yc��-9���9�����[�U�a�.FQp�k3���
t&�Ey/�x���o��jf&�>�W���P�{Vhʇ?�z����=K�C�qW_� �7L�@��9�K�`�J���y��྆�OE��3A"��ӂ�|Oq���z=�Bn�̲�nv2��%�אu4J�$��-{RMХ�c�x�����uwhYڀ��i�MM�
s]p������k��G��}���,����n�	�o
�1Vl�+
e����Y@^4=�k3Nu�υL$XO ح෥Q}�\W��u=~�V�E��G��(�̞�7&m�=a�p�����X !������s��`E&G����<	1P/�x�<��Ť]���*]��� ��X��	$W��m��a�U`ӈ����������H�贤��H5R0��$�h�e��4��8t�=�Sd�DB�[0r��
/#̦� ��ŋԉ�k:F�^�����;ݮ$��YQ]�M�"��P�T��N�܍0}�R���Xp�vQ����ѻ��?��l@�std���J_���"ٚS9�`�����n�2�?(E���vf��'q�&|���d��psO���'(+.���H�B�Y��#���Pe{�R'��
�[,q Cw���{E���J=@Aeg��p��vc�C�[�WoEw�0x8�G1a7yg��)S���A�=Y�`������M���s�}���D�Z}��&#� D�v��ʒ}����Uݮ�v���4<�� ud9胥u�F��G��|�a4Y��ĠЈ�%�q��D����,�B�܀��@��Y�c����6�x� ��B�t�iN�ۻ]~@��g��:���tY�'i�	Y^c�ua�J�d�-���ρ0��
&Iip.g�3g�O���+�`F_�!M�C+��-��0���m]��G��j�JW��]��ǚ͑�c
�Q�2��ˌ�Y�S���CK6忳>Jl�D�)W0%"���#���j.�T@���G,��^�oz$'& ��4'o�s�3ܶ����6��aT=�H�l�yC{�(rj7GEJ]L��o��U�W�}F�O�rC��I��@#DI&��%�~�P�T���������!�A��;]��8���p7̦�[R|D�3]}�F�ԃ�+������]a{���P������f_�s�h�tJ���W�����"^iw94�����~�Xx���U�pi�	�8�/���/{!?�q'�H���ߞ���	�g�Y#��ۛ*�({���:�巅(���7]~�ClzO�co�_���s����������!n�"��6�Uu�J8�H�1B�O`���4�U|����$c,�����5�Ô��Ȳ�#s�[�ޝ�2��b�b�Kg���j�&\a(����P�I���(DQ\m �� ���_��g��b��ia�+N��M�Zg���d�����' j�����&i
cqx���+��=2U9�|�^ܭ[��XK�99L�*�u�0��Fd��r������S���&�bf����{�v!婠�0��H���R_.�՚]�b|jǢ,��(���F�a�ջ2+#�S4&6�J+�)a�?i��o�-��ÿ���f����k�^�x(���ak�,����1i�����u��8(\�6i`�I	/?�����Y9���ݱ��&o��p�m#�4u�,Z�9���8������|5�^�A~�8Y��J\(�j�9���r�?�M�])2%5����K�!Q�ӎ�L�	�9�g>��\o=���m:,����hknD	�W��N2�� F�;�x"�s���;�rz[�h]��^B��*&�/�����hBGBO�#�&fEtQ�`;a�Ӥ���p�G���h����QE�U�)\`c�+����,h#�S�Q5�THAp~bh.�˒h�AdvX�v*o1�/��}��`ny�#���ĩv�1��K{#�R�(��O������+���ҩ�����x�
Iv@�}&�M2v�Ps��x&��^�p�����7CÉ�˻������g��A��|E��U�_��y�K��֥� �yr A����+����P�?��O�;{Kwk�qa�Rnx�=yD�lP���+"M����yWCA���Ƹ챸���L�����ni�����L^�"�l���u�Li2���{���Le�e��Z}k瑁9�@��/SC�d��xNwT�1��9�v�D�����%����ʓ�|~?d� ��0eL�hlue"ߨ|���O�����:��H�F�!Y�й0o���.��
�R �d�´����4Y�"�~˼�Z���eQ���������� 6���b!��o,x�Wdu�ݵ9����`, �p^c)B��ʃ���nikN��s���/Co=�*�=�W��&k@��8��Q_(�Ԑ����!{�%ok�o7/p��U%f�^��O�(۷�D��Ʃ���o'�?yD*:�A��ޤ��4A��:�����x���B!RM�v�ܻ������t4�	�̄τR�袔�fg7�v����M-ˌn�(u��7 ���8���s+�2��I�Sfl@.�Ww��-R���-r �ɖ����o��@�e���D�#��~Ѻ9���E���o��!�M�X(�c������v��;��u� #efW�x%��g�(�����8��nk�>�8�f,��YԜ_��#��{���x�`y���,�k��5����
��t�	+lȂ=
WbPÉ
�I���l�u���,�"���a"���[����٬��83E���}c�i�_W����K��(8��[AA�VpY(�_c8��윥$�~ᇭ+���W����"��]t��y�-^�`��<�p�n������E �}9�|2��˟����G5g��$GF�w�kKs`�l�`���
�0Dj]�Χc��6��#�7�|���&yf�}V�9����!�xzU�t���.�%E+���H��9n+���8_-;G�#���	¦�)^�S/�ҧ��jmg�G^f�F�%|g��ݔ񜏠�,�I�-��<E��$��i�@�p^�H?�h��$������!�_,�i4�@:` �ݺU��n�	YCmE@Lc�� �������尼Q�9�
]Nk��&b��
mHлf=�f���,������\��5��fC��o�W��<�-���������St��,.[���7���=w��!��z��������c��'aH`�����:rEn@aՕ�P�ǐ��-iá03��*�]�ZHSN�����@��V*P�e�B:�
��[_x���F&y���
�w��+pe����!Q�aݒww�i���2]m�a(>�ioJ]��/O��.��ZO���gE�w
!����Lx��\��vU䢱�eg�Ҁ�k���pH����F>5wuTl�,�%*�9����į��s��I*E�����O��;�l�)&���0zZ�����ǩk���� <(�8J�+|�H��zA���J#����0��/�� �����BO�\���(��5M�#Rn���G��]?����?݈`ؿ����yv���k�$������P1ϱ���e�؛�E�u�@�_��(BL����L ��h�t�Ko�ɳ�/�	(7"��2׳�Z���Fe1���o��v3���zs0��dJ_-�Y���P�sS���Ôh7��e�����pP5Oƌ�OB���:?���^��"{�V�S�I���#B��ޭG����_�9�5��_?jy��(<� ���m��o>��O����d2�!��w{2��5�u��~��3�Z�L�R���
�W���U���9�'�nٜ+C��1p�)	׳N��[IV�:��e��;�r�"<�ƺ���%a�7���E�kQ.f�����:ָ M�_h��a���C��z^���#����F}��/�*���b�P�ga��O8[A�GH �w��|8��!!k����l6��&ܰm*<�VV�8�0��6$�NX�-"�C�=A0g�s�������O:�K��>�6��OQ2�om�]��y����$��n&���4=1P�X酊��t�Rt�/���8s'�.� �g�R�8
��V0l_F�,^�{]�Yz:�L���^�p���Y��>��ߌ
Ph�m�u}̽v�ɜx}g	ww�!WU�XBWeK�?�>Q{�2�@GOj9�^?&�u����V��9���B^������k�9z,�2�(;��Y����|�	>V(c���N�&L]L}���F^,��N���M�U�G���ȴ_#l�}8/"���#�GְP��1�6+����&ò�Pt%�RR�}�\��q��j��ndK�-��Cȼ�y����z �0�2y�7��d��{`�l/z��.�E��Gv�8d�TPRE*A�E�!E{�2�_�Ee�b
{����� �!u`�e'�Jk��i�yO���4ߞY}]�� �{0wJ���K�t�0޷+H!�Hu���ăB�kL�@��"h�������v!S/�G頎4
�v��n|J1�'c�Q�1�Ԫ[��q��emq<����K���M|hѼ�A_��+e
�WEO��[/C32s�j7k���D��2U+J�e.�	�Rk�dDZ����]��e�l�7�� �v�(��ؐ~9hCG�)	���{��V8FaxϸL� ̃<�D�����	�rz_�� .Y-��j����NЊ����2ŭ�QqY�Iih���5;��M�G��	3Ķϊw�t>�s���S�gj`��9g�~�;�/��BmB�c���kJ�V����Q�Б+�&�y�!6U)��'�{��s-*��|�Q�,d1�2��d��O�P���8-'�ŰЋ ���j���Y��~�t/�0���it��Q]�/NgI�jV�M�.���߿'��PT���U	h�'
,ȋ��*K�gF���؛!�'jJ���(;"����YCk �� F��6?��ۓUN�y/�����E���0;�藌K��,��<`PYP:y����������Ј����3��n�^��xE������g5�~bF�N�Kg�jgw�39x�D�?+H2�4c u</ֶJEm�x���p��Y9@v����*��Á&�$���uե�U�,N�l�wGMĬ�T��e&/��)��JdJ��?4���n��2J�u/�8(E���t�`�h�_�D��|c�R,f"�f�����	��$X�B&�����.��G���n�Y����s)#�t�{;����L�2�x�U��V"��RW�B��a�8��y:)� ر��c$=~��a~wC=�]��:.Y՞{����Ġ�j*�	߂����xY��\P���}�39�Z�%g��f��HN	��L��2/�T�׹�8���-��B�azw���`��[�mb�*V���G�m�&".�ա!Ԉ��1o'�?��>��H��o��K����>�J݆ᥱ;�PV93	=a���u��<n0�/�Ċ�7ߋ�FF�|�L2����n�P��;�&�E�e[L�N�[?���U 9��퀅i��LG���ͱq �4�zVi������m}z��u�9�ј$%�<B(`�y�ޖ�t�u,�<{>S)�A�!b�ʅ�Tw��5��"�S�����HJķ���\����=U�:�l)�haR4��~@�L��N��b�U.-
Y���@��P�V����:8lC�W�8����DԨ5浲+�f|j��W0��W��M~��?zx��lh^�Jn���\��f!\X�bsr��H�������=��C�wE;���n���X7G@��NLD���/:~�����f��IM74��k���5==g��r��~�w~9�55U���u#����v_.ώ���������=o�f�@uT.��f�����Eg4a����T�+}�ߒ��4��e:H1����F�h�#��O�t@g���l��P���r��V��99���lw�>�&;J:�M9���<lj>`�� 7�a^[�u)[�.z�0UM)�s��ӵ5� d'�C�^��蔞,S`AP��Z	�Q�MS���D.��߽,�avrq�c2�K�d����ӎs��?i8L���5_���~���{>�0�~��:8����w�EFj�/|��ϟ��_G�����-y67����:T�� W� �o�����ClvX�@�-���$X>�+"�lK�G�5�O{d��a%�xH�Pl�"� ��r� �b�YQj�����y����cW�~�mJ��?���kF���2��i�Ǹ�1ؔ�O5�'&D��%J�;b�V��~��/�=�5~���ݠl?<�{���4[P�%e���A
������HV�H1.]�*�q�3��@~��X])l����!��f����Lg��dd��\[���������^	:䤖ضB�S�PE����c�Q�8x����t�y7]�A��h�]��?��`�vG������J�m9�-��6�f3Ft-��S]L#��&{����-����׍F� `��?y��"'�*�A2�)��j�#��ņ\��%��Woly8,q���%���_�Q�����VT���c"�eĞ=ؓ�z:D��$���P]W�a�<����ү謇�S���`r�?�N��otXZ�G8;i��(Y�)�2���_��E�Y���aMW��^��xk��y~��O���ԍ���:Uҁ�03�ٕ���lQ+g:�;��fϷ�%��#���! K�8���e�׈S'�N=�����@59�f�EU�?"�Q"�W��B�m��������lXR]g�ʃ�Q.�_�\O1�\��z��I�(�	���he�Nb�}O	{�I��j��Pwd��t�}�#���&�@1�'�1��=���x�����8�`��S8�컩Z�/a�X��N�Ƈ��4.aDf<H~��v�}��K=�������+����u�KKn��=O��Y,TJq�Z5�R�}יF��o���{@���M4�^��O2h�(� ��M�3�@���2H��5��^�}�b�^��@��O�k�Ĥ�[�e0&��h���T�ǰw��A�g��L��J�n#�Ȓ�c��\�+�c�j�v�Һ�^B�b�"�n�e��֥� �y��l�:�s�dې�F{��־��m�O�[��5L��c���^������z�MZ�����k:���!4VCQl@	Dpo����벫n�M�Q�$v�ǰ>�{�������/��n����ey�����p	Et���,	b�*`υd0?�9�1�}%R ��\����&��xs��=�W���	]�J�u�\�J=��,C2,`�)�[�\����&����ML��,Y���j�W���v�zD拉{Ms�AٺVQA��~�5�R��a����'�@�iף�q���]��E�p�v
�4�jpW� @�+�l��b�D�v�~:���V͔v�茜�� ��r��u�^r�r�&6�j:����XOoh��)D��#�S��S�:*$��"�o/Ͳ�+s:�}�J�" Q�fP��lU1���T���!�f"~Q�P��)�$N3����5+�=�f�Yj3���n�D3�hMk���9?�F�X�I�{�ja��Lx�`5=���g/OyK&��O@ }��/3��a,����"J���=�G?=hZup*ޅT��5L�y�$���,�/�4�n��tI5��׮V���J�@h��bY��\�B
!�X֓��M�ڠ���+q?ݺZ����z(��`%Z8��dg��2^R_8*tvoD��Tғp�
������B�(�/���h�E�^Aΰ��/�>Jz�M��k_��6,WF�
�*R��
�6�(�m쇹��M�c�N �����q�u���L.��j�Y���,J�M�1�[ߠ�3]�̐	�NV}v�#�V�	}&�G����Kd?{V��B��+���@'��6eNXMjҁ����}��%Q+Y�h{���(�'��ӭ����b�\�ߵ��Q3�~��=�&x܇�� 	�x�A�}��$�uu�_h���
�1`�=�x��'�{�����I���v�@��l#뷙7V�-�TJ�
�Y[@�V��-Ej|�|W^#raʘ�0�[�Q�7L��(��d*���hR��u
���U�M�T����Ft����]|���CMA�T$هf�_,)�q5+���I���{c�l�� �*���xB%{�����YGj�J�w�Ai�U{�}��SL�<ssz-mK�[=|?��3�4+�Sv�?.(u/ �]y�!+��X�n�V�sT�������sVr�	ʩ9�q��.d��T��Y���A������]�j��q�2��z���z��F��#���9ޭ��-cқ��]-)�鈎ē��HU�`M\��K�4R䮌*����)���;:>f�o��˛ya�U��X�L�K���˜�4�4gl�\4��M���(ۚ���KP�	�M ��8X���ZWSd�&v�.�n�*��tm�H�y��ZrP�H2^<+.z�{j�'#:� ��%P�9����N���ZI�+��<�.� 1�x�0�hG-Z�q����'���=P�c�\�$uF��/x�?.OI� ���1p˿�4��&��C���:� �<�U��0Kv�`��c��[YJ�5����\jR����Fޱ��~m9"e��ogX�T��#m�8w����Q����p����R�-�9�,��ʣP��<*Т��%��	Jr��>W������)�S�=�'Do�KM�R}_��=i
�0K8-7��*w>|����b���s�#=�k��w]�C�`+�������|H2�����Ф��#�Sۊ�\����c���~Z���zp�ч��Q�YjF�jܔhs���p�*���^
�Lo����3�.wx�����B�	���zj���+#X��i��~ҷ�4���LF�m��@rI����U�YE�Y��=+�-7����	��������eN�Τ�I��*F���YU�/����TF�IWOXS�{���!5._ba�L�M��A�y�q��>	��.s���WP/��I_T �
�D�i:��=W�ѵ�M�dt���ܒ�<|�u�J�Ǜ�G��A�Fa변 �p0�\�/�Vdқ�3.5���8�K�Di_��q�n맭���x�'�h�90V��K_)��!�ڨ�[C�t�w\���@bm9X��\f�h��'��
VM����i?R��v�k�����ImR&����Ţ�o��*��׼M�H�ktb��+�,3ҙY�m���V0ޅ&������5O��fI����T5V���;�T�<�;љY+K%�K��> �-Ǡ���B=j��P��~Nbf�ӓn��z�̜�b�3��G�m�"�֪q�y#<�^N]�`�~?����7��}9�D�*�X��N(��ď>��r5�<�^ꛀu|�T���]9��n+���!�1�3��Bi�*oW뚈����ڝ���U����h�Tjh�tl���>0K��+qNrvS�����I�5o/Њ~F��
�{��2p�+E�s��"���/fnS<<��47n�l?��,RU�Hh�r3!*�}�GA��KY�: B"�}ΥA�1�k��);�!L�mp|� ���ߵ;1B?y���l=�)�e��?,3䟭@�{)�l�k�����V�We`o�v��h\كc� T�M�@��PJB�@d�GVAX*�Y�2�Uf.�a�Q�:нL&Ϳ՝/����S���eK$p�pc�עHŌF��b�ѫEd�?��zh�9}��]�&��p��^�����	�o8���ʗ9�gT-�83���C�'r��ԁ��� ��(��Y�����.N�Y��$ҭ�ʨܖRp-�9��� �cy���W;���b���e��B0sÈ��L����sH��1�B���`ى�>����1���;w�t�]�5����&�(U�x�H���s8R��Wv�t�����M�Β�n	v	���b�~O��P*ipz�ٍ� g�6l��ļ�w���-�*���FXM��YO�h��EnQ>#[�����GS%y����#l���t��e8���� Q�4E��@��(��� �α���i�m�������N�DV��H�/���Q��ey�̍�'օۿ�s����4.�B��1�p��
H1�������4�����s7��J{_��i�"(G�����iu���7��[�pǦ�Ղ�A�7�T�3@ ���1�5u��BS����sNX T���yMgHW�
��_$���c�D}CؤQ����Xwa�'Q�1�ҩ��g@�墳-���2�Q��	�H��8��lĕ�X!M�����t�g��i�=8�5L/~�\޳��J5y��X(���k��3(ܑ��E�XtD�$PL���]]��CDƸ?���vO�6�I���R��iZREo/�ښ�Gm��=��w�m�\�w![�`V�����eb`\S�,�|:���P)C���D��7��
���ր�U�]���ȹ"T�O`iA�@�w������;<}�������ʋ�9�b��fj2 8���$��A$��=����ɘ�(?[�	�H���=����|�DEϭ����#��N�[�Q�W�AM�K�Wl�4�G�n+�g��e|�vX0c�e'�]��ƍzf�wtY5F�՜ME���`�6����\����r���b���.��g�t����do��`\��[s�\�I��`����k鿉d�?hM\T*�{���ː7�x����������U��x�U2���K��hO,)#kD�D����(�����*�Q�s����r�%����(���hP/%əC�-�-"=��������7C��=�Xd��On
�<���� �gƖbK���e�W�j78l�v��EB��P�Bv*�	һ5�~t��w�霫�]���Q��������<�M��
"!�_ʏ����n������1%¶����IWT�2< �ëK��/�h^�����qj0<T+�c?��/�����-:�ߟ�L+�ZU	aB;�[:������+����5	���9iD�VIt{� �>�u��|ap��.�zW-�e�`Bk^�p-��`i�-�,�������^��֏�;q�q���\w�@8��c��p!�"~��V��>Na`~OCkO�7�:w�l����d�Ǐ�q?]���#F%�齇H�\��[4���R�xyv,�3�#���$�J��cEH5����B���ǲ�����"��S�}��߅^F�s�8�:A>�}����ٟ��"���>��\��� ���=_XS�ew�4Y�u��6��7�A`�E�1xg�K�~��0�"���!��0o{Ժ==�����6���+ڬ�]fh<������bi�C�����w�^��2��mO�Sy��q������ ��zh���=��e�_5�2]��%���О���^���Kx�(�#4�)^��Vv�g�`߈�m[�Wv�1�g�m��sJ�
���$�v�Ig�Aa���YV�~k����$��;��~O|�Uӄh��Gc�.�-&_��OJ��\Q��G���I�A܀.��衻O�����0ʻ(�N�!g#]�LCֈ���rq��fi�=f6�N��/-�K�[��5���0�Ã:D᝺�ق����\lƀO������쭣�
fX�'[k;T�ɞ�ZiV�r+�n��|��쓸��?axr�,2��L����.Y$=�?��-4�̉B9Zy�	����^yoZ[|�[:�j��{#����F����w��9+����A^��qK��D.��}�#W�!�?E%�*�.�l�A�]�'T�O�vQ�9��m6�N5��ݣ7�K�>z���Dh� D��>Rэ�6�nJ8�MeyF���3�����`����z����+2��� 4Şa���;_I��5�]�M��6XV��-O�ڬ'��^R:��)AU�:�v�O�\�+� a0m�h�����˰h�(�-��E�ѓ��#�F?;����<>ttw�0Sѥ��xK��Z��πzM����IHg'l���=9�q\����g^�����m6|<�^̛��16�_�����4y~ɼ���5�����_��=��%�O]��4�#�Wh�0��,��GV2|R�QHA�]���\����J�q��*�z�������%lT���-tJ���#����5 �C�ܣ��	�hO�	N�������i�8>��Y��Q�ڎ��^�㚂���	� r���Ѽ�ET��6��8�����HqV2�@qI��Z'��Z*�i`�$T�SG�̀h�V�w��";�  FZ!��{N�����e�o*��z/�1�0�,�?=���{\lV��H��`��%�� ~ۢ��W��c+t�4 W`�h\�Y�&`�+����3������]=��uR��j	nd+Y��~���*�c���M�{�ְ��n��{:���T�s�:վ����L�LC�@��K�d����%b�.D:�r�,�G�`k4��ҽ7U7����ƶ��G$�U+h��wVai��q���Pds��Kҩ	���sB���
��q�9�:lʀPnE�E��&w���Z�ҁK�JEQ�,�V9�72�"'�ӑ}{�*�IƯ
���/9�O��ZY���埁�6R֞���v��Ȧ?�$-6���	^J�h"������n�V����9��vD��scR	�b�;VK�:���xv���X5��r���Ɇܧ!π0^�0��T!�I�X�a�~7�!��L��>�ʕp�h���q�x�1�~����-�����vB��]�p�l�G��T�jN��f�6��v!���Q�*�d���3�l���S�~o��7�dӪ���u_����\�9 Kw�fM�[T�w�/��t�(OM��J�-CuwzG��G	���4���Ǹ�_���TM�)S���HLQs���s����$��'��PCqÇ���h��8��5�0�A�[�*�Һ��֢�{&߫z��&&�i��n/�J�W���ru� �����h�2iP
JJ���l��Ӻ
{��x�k��.ڀ�����E�:q'�$t��y�JG���Y�(RG�D��R�[
�j0gKO�j�6��Bp)u`�M��^Ǚ#�O�?���e!��i��
n~�k:��:�/���4������ƾ~�Mx��c���=�ЀrK������qi�����R-0��J;�o/�K�/) ��[:�Qwr�[��F�K4�vG�	��s�1/y-�X9�kR�2[�Q�E�|�1��b��
i7��U����1pE�;����k�t�Lb(fae~n���L2a?Mࣘ�a��{�����y��"��j��H�=�7��vV��c�l\x�r��F{7���z#HA)�!J-�1������@���<P�,�����,�|WK�#J���骲�TI<0��������%���C�^�3�)�'�jm� m�����e�b"١��v��$;����+p�:�7�� �9],m�G�����0pS���gM!<k܉#5̕WD�P8[��i�'h~���DhÙ��d��ޱy�$V$`.��Ķ�eO�ꍑ�F�J�(97�xӡ�;1x#L2I���)�OM�r�����t�����#�D"d"u�xJ@e�==�\���2�K3�-���"]O�����=�WV5�F�&T_���8����W��,�i'*\�שx��Ш�@�ֻ(��$Х����u$I�R�<�A7�l
G�����n���d��iHV
��O����� �sm
��B��Q���a���;�c��d�"hn�1ː}�Z�Z�S��P-��v^1J�(�t�_�{w�z�X�ئ�&�.��s�R���0���u���P0�/�H���:�ﮪsw�=�~������:�����+:�Uq���,u��
ۿH��:��&�[)�z�h��мUV�뚎�T��ą��ϡ[b���f]�KZ��
%s˹�G���Lm5�M�S޹/%4*K/e�'�����#�M�:l�XA�����W��������j��B�� �(����NK�T��x+k,��jA�N1K~��F��0���k���i�)�cv9�`�r�"�~�5WP�M����f����!�E6u6�|C8��-'�HSP3ʨ��r�m2 7��m�����5_�[<��elc̜ܬ�̀?k���&ƈ'����y9;���~����@��X-�}�J�[��E��
�^Z�X"�뽬���I]�ѩ�o��t�`��Y�����l<1c�.:��ݟ�?��W�n |����r�(�g.��+a��>v6`ˀHp�^� E9�2m��lB���:6K���%Ep߃�[5�*VQ�g*z��UVq,F��?��hgcb4uC�����ғ�_O�2�7���#��r\QZ~e�S�Q1�Ł�q�K������H����s N�P�x/�ߵe�������?<Z/�~KQ��yM]E{�hى����m�����2���[$]�攞����+��xE�^��
�4�u�[w��DBh�L2O�>�Z�C�PM`��y{�/�M0C�m�j��x�P����ʘ�d{�_����;1��3HC@\���YzW�A	"�QjyƋ����g��%��@�w�,���W�+�f��3Ő�.B�I�l�W��?Wrb���He�}mn�,e�ԇ��}�j��CJ�;v-�k'c#%B��d���$fxi4<�/�V�Y%���9ujy'�"�q�\d;d9�}W�ξ���R����)�{�� ?��ӏ���L��eِ�a"Z�S���Y��C}�,&{ǃq���Ǫ�@u;
�i�C|
V}q�һ��}�gx'	~��֎���\%P�t!�~Y� �N���n��:15�`C4���SK}��5��۱��s+�eĐ8,�Z��>���^�y�`�^��K	�L�d��8�|1�1�x�qThP���Ɵi�#I,� ۿ
An�w���I � ��6�����(P����N��u�]��n���Ƿ&/���l�uҮ��ܿI��J8&���!���&?�e,rz!ޚb�V�&��Sx� :�$�l���}j&�x?	ԗ6��p�Bl���x�Flrş*@G�l�H~A��A<��8�Y����PY;򡐘j����h�<�}��^�5�B�����sGL'���9N��[���H"���a�o,�k.�YӤ)X���4��<���4�K�q���C9L	՛�L�*յC:4j���ϩ�xZ�<e��tsmz�M`p�O��l�C��Ȱ�u�^ַ�~x��E��O��y"d�W[r�nԱ|i��T��me��R=C�Hڑ��ϐ���3g���i� �BN�Q�;!�.
\
�E"o��iv^Ü����0�C����9kb1���0��#�`f�O
��h��+󠟒ߧ�w���In��<���_�r�i!��&�&ۈ�b"��B�Bx5zl�����L�z	:�*��J��Xo�RA���R�.M�]�e��?�t�%1�	�:b�&�h^<��M�Hz��q��ᗑ��4c�AR�����-=~o���\N���{M����r)I��!u^A���|�0#��Ų7��b�V��]z�[Zg��% )~I}���q�r�J9���G��4�ȱ�m��[*�|{/J8���.�-�F�H)Y�datB�Ed[^�"FjNh�0�~�e�D��Lɛ�v��w������`[�� :��r�U���1Z��Q�<���5��wi�E]�3ҡ��~e�I���P���x���S�ۧ5eT�}��č��tB��MWO���gWd?�����K��*����Wv]5��ؔ�����q*��
?҉!���D�v^S��16!������	��AO�P�Tx�*d߰����9�uf��-���&�\#�Y��.
O�!G�����~�35��3r1���d�o��@����� ��N��[ڎrA�K$�}6�p+�5�౿C�Ʊ�ۻ?r98��_�6���R�����"� �2���|T���*�t;�!�n��>)�K��?��e:�&�Th�"���x)n�Tj�݉5q�=�[␑����h�_�1"��.0،�]p$��2���P���^��|��u(��߷�@0e��0(�^�o���B�:�}z�A���a��[�<D@��H�	�o���s�5�b۽*�7-W0&��%_���q�TǮ@�K9�M�n|�<�E�b���(<bi5��$>��7�`{)R�۱���᮫��UY��fJ͉��rm������gf��
eF'�Z�qpC-ogK�����6G,�{+�ҿ]�7�XZt� yM;L����)oOv�zqI����%:�����}��۩��;]N�f�_�� >5��u��ĳ�g��#�����g_G�$���0��#*Ѱ�h]F$w�֩o��D�ZJR��N��;Rq!���Z  �w��.A.7<�!�<��C��\�h��������������˼�R0�M/E5�˘A���U^m㼠�U��&�7łIM���>6Z���������<�>���6z�R����DHaGpy��-Dl�:Q6�L��8���ݔ�vE>�h�L�]�S!��!��(?g�J=��j?��� ��]�N�\��5��wH%	�����uk�\�I-"7
y�!�H�p��JGBu�Ӻ��Z�(��EݵE}'{��=ҵ�	�%2���Ҵى|���?�y��2�3����H�W�Y��m��)��ŧ�Uk������z�[�׎Ԫ��#�c�$�U��9n���n�k�KҊ�ܸ��5�5.�����f7���l���:?�7&o#@��*��bF^�E��|�N6q�]���n������*6���l2��^\hZ]�m�F�N�8e����r�`g!��n
��+�;�G(�[�$A�>�e������^���;�|�D�@�GT={i+��S2D%O��I=}�k�
��>�|���uD�\sJ�Տpˮ#>�t��Q�ߖ���v�qm�����W��n�9Й(����#��B�,�Z����2�>r�H�<2��m��'�%$QŰ�	���/���o8
X���������d�k�<}�ϸ�ϫ���B��]�� ړ�(n���1�S�Ή��f[�?&(�yد�^�w�8�$��>��A��ݢ��b�)�^�}.��oV.��bL���9��^�$���J��齼�}�8�eI���ȿt�wH⚈u��n�إ�3Fn��E ���]�iT+k�P?����r��j��%���N$�"��k���[Gop�
�(sؚ��9��;�yn5\{܈��5P����{�Xz+����+�Xm�~�m�p�Q�ɕU�bD���<��� ⎘{(7�8�)G��&�d���������,�鏈�\ո[@S������yx�|�A܊���;��­4݇Q���ྵa�x�D̏"J�$r�j����u��FM�vhzv���F�рn��Z�m�R%���h����L���� 1�`!:p�Ne�̞�	�t���S:��E�zHgv�7c(������7o8�cY�;�ja���r`�3��;�G`��U�P�u��F�1�(�{~�̈́, C��$R�����g�`ith�]X��M�%9�8�P���.4u��x� �-MӾʯ獪����V�+�(vʛw}���}�+Ӳ��5����|�]�������v�?
R�ܗ*{����5;���������!<X�ʨ /�7���12��h
ƼDY)�� <K�Y��0��䕋��dъ��G#c���Uf��Q|.t�ȍ�ڏ���	�q��lq�F،���<=��9�+�4<��/'�������*�>��H`�?D�f��
Sb���Am���ِ���}�L��>Z�t���W�ʻ�,qKOO��!y_j/�U,]���n}:X?�� Iڄ 0�+�WdU?ҹb,���46��Z�>��"�j��@��"F�%�bxUm�`E"T�-��&6�o�Y�x��*F�b����Ґ��ا�d�D|��8�ܚ��d\����Gt4�Ir���[���sD��� ��f4Z�]Zr���(�j�	P�CV��L�[�q%Ӎ8�*�|���)-g~.b�k�j�j��V�VHڂL#J�r:
N��举�1�����R�.\��i���tTn����8�d������Ed0'��R[O.�8��F�U_��&9O���m�l���d߁h�1s�g�Pj���y_��kX���N����b��S��� Ā��.�:dB����J|�O�a�G�����l��^I؍##ҳ��h��ı����M"�{��Hs�6��1;���TT�e�EB�k�^%\�w�ހ�ā�e�r����U�7�u��]���n��5����6��/�wx�5�u�_�B�d�Q�8\���=�X��鯁X0ҽN�!ˁ9���+b�����$��ງ��o�a���|0yvY���Kt|����epIqZ^�5�1�n!w:��	<�z㾳��(Aؠ����I�w=|�7_kt:�`�x��7r��ȁ��t۱,����Y:����zP��{�_���HfrK)�3����Ɓi��]*m�yT8|'
�-z�a�k:7�l�_() yy��% � /�Y�iVH�d��oH�*�v��z��Op[	�\u�uM|I������إ#�	�U����g�c��>��s�cFm���~��s��Յ�\��2uٕuqO������p����*��Ѯf4խ:��ݒ��ō��>��g��n,̻����v3�JP�NQ@�x1.���"R����uP@���U5*�Jd���J[�䓖Z�ϟ�{��I8S�6Ʉi��ڼ�O`ѝ������Cf�߽���
�3����zV�����
AeVG��\�Z����Ef�4���)��H��ҷ�T�h�cT{�ug[��#���O�f����rvˎ���>��D{Ͷ�թ�X�kvK��,�,��LQ.�j�"K�ߩ�ܫsi�N�L����TeT��ծ��N���$}@�<1�xb0p��� ��vS�{^��}���q�BQ���N��ݳk���4����Z�u
���� ���HH�Ϝ��=��|���=J����U�f}�dQ$L`�C���Ť�A�B=�a��~�@�I	�͝Zk���+?	�8wp,q���X�Ͻ��@?rt���p�;U��	
>��q�̚1���|�����^�%l���r��F�"N�nY�	6Hԁ�j����3�V4���R�^����%��׳�4����?���ε���������N嚚p:�D�vc���=�����ɦ���x��}�+7�
I�H�P6���3��/b$���EZu
%�
E ��~f���ݩ�Ǯ�^�Y�3�G#"]�3<�X�̾���������zu��7O�~W��nGW�.������xx�50bjn�d8�{�멟=�7c��*@�Ev�Eƫ�&N�T��.zk�Ro��u�l��x���Ll�I��.�c�د$F8�����`i%&9��(���NXRzj�ޟ��)w8bP��}�� �j����b��x������������`
;jԏ�zvm�`�Ț6?�O`6����#��b �!c@��&��%�:�w��"�gE����Di5�6�|PF�| �?��dd6��{ޜ��.ܿGS	�/����PoO亲�|ٙ�>�|��2i)���hQ����@�E4B�����V��&$X���NL;��d\��{@��H�M�d?d��]���4�qKb �8ء�w�}Ի�X�7��
�Y�c�mr�`��m&��j����њh^@��v��Y�*��
�԰\X��cC_�]8s�N:n�T�X��<���t8�j&���G��<W�仍��
�lq��������E����L�n��(ݿHx"*ʭ�������	��o������u���0g��Y%�>�S�˜)ϖF"��� �/�Qs~6�2g�2��l��	�"��Q� ��
�v��a�%��\S��a�澯�r�k� ��a��w��Ķ�,����Z��r8v�p�p)�%�@����?��O���U��ɗ�ƛ�D��S����?ȑ�=�c(P�^۹��4�#�XRUD��B�I[\FxޖM�~��%!"0�:��	FAء@����d�u"��}	��\@�̈́�5Q6T��)4�;Z�
=K࿟��y���t<S麽t�+����
���u\�����;�j�0
ceR�QxEq!AMsY�b�9 �U'�)Ya�,�[�c��\��[���8C-��pJ�M_�������c1R8oL�`���^͛-e�"
�/g�n�=؊�=���y5��4�	�
����د��O�ߝ�x���>���#�l�6W��?ird���U����[Ґn��[�褐�q�>��L����i�ŋ�a�3K�ł̘޾m���b���)|�?��Þ����M��=8�.U��s��M&�p:<�ϱ���՗~�hW�����m;�&G&��L���w�����0�`3ޠ�ݱp�C��jJ²
���Ys~�2�k�-�)�,FX����P0��5R��SP�9�I�d�y�~���j-լ��t��h��*�&Cg'E�,����w�A�T�#�����?�|.�k|rY�=P�B���S9h?��S���b]�?��h��N0rw��~ܿ���ͣ�Z��W:��_�r=PA�8Vq��}OԦ��ݿ8θ�Q��lCN@^��ܻ�g?:���@����v\B��䰦��?�r�L֟���@���Æp��vS��v�N�߽(zC?��-��	�n��z[^
�7WT�q����r+\&�A��	@���ֱ�sg�2���},�wu�9�c�tP���ݢh>#�*d����h�8a�#@��a.П�g�F�6���]�����YI��~�Ȏ#�E�v�crsf����� ���̉ ��a�������j���6�cK_�.!��pJǁ�AW-�X��+��*x61
���"jC��Z>?Y߳W!���$�_nK���IE\�|p��i�ո��}i_>:�[�E���	�aL�F>�
eZ+���ZZm�����q���؁��jÕ�jN��.�Յڽt;�B��Iq���3�jY*qW�8P���I+��)�p_�;��EㄻO�G�@�-3���?2�*��1�EPF��mGc�X�'�{���9?I�'����H��Ƒ�w,�m�fr�Ck���"�)6��޷�G��gw^�x⹡���v��lGcV��~r�njaK�o�V�g�v\nZ��ݷ"G�@‎y/|�f6;|JLE�l�J-��]��Ȼ(S<� ��ѭ(����?� T��
�O�9`�}B�N�rU�$�(�tj����&e�!�Q��57e+�q蒢����_�B��T<�.8�O��r��d4Lb?���@k(2>G��J�����f���?��.
iA�Bf,��?^�'�(3V�m�%�&�K�/�����<����l���IMo��~���K����g��#ý)��	�e��Ч�s���:0�vkWm�G�z������ʏ؋,Ֆ@T�C��|�8��dQQt+�.'{�.O��8�ro@��0/���� ɫu��@Lz�*���(����[�Rkqo��*� �lG+I�Nq;a��6���m��t�nX=����D6pwFQ$�Cx����g�F��K��a>���{58&�<��J����| ���Ϝ�W�+�tAE��Ǐ����t<��3������L��mh�cq3�2��]��,�ƭmz�tL=M)a��f�J��%�"!a�?�ۃ77r��k��o��d�a�Ӓ�����`�g5���f�� �r�M�ײ7�m0 �ʍoet�`F���6�'�c����
����e1!� u]P��-�Nw!��y�����$މ\C�F�3dq�Y̑���.�m�
.�B߼�E��$�ϛ��@0'N}���0yC��CX�k�ma3�dٚ�{t �4�zR��Z�y�jV�������>c?����<ue���p�kO�	)��dǫ�.�����CS[Ԩ1<y`�+��"-���[�ۃ$� \�7��v�.�������1�Wd%�^��*�7� �TT������ֆ�փ`�D�iO���,�3˾���OJq��[��+�oZ,��/� k�z�y���D�����P��o�\f4?��h��_"�K
��8�&YUƢy�dL%��7Q��H��˓����i��L���~�F�Z����L�~E���1���Y�R$@��'k�wFJʐ��y��ecǅ�A�G�(+`�?����+(q'"n�	-qю���ֵIZ�������Knw0�b ��O�Cb��'����$*��H��� �	 �B�SAu���#p?_��T��h�fF��,{�t$"Li�T�?L�E�_��*
������2S��<d���]Y�^"�����h)c�fG�&(��E�]x���g�� ��ݍ�]�\��m� ����A+�Ү�
pMm���Y�ʬ:����mQVy�:����yv4���#�8
��1��+��a�:�<-� gyF�E�����V;�H E������ wGZ	ey9u�Z��o�e,���c��贫�V�W��8:��"� ;U�c�Ա�6��2�+M>C0���0��3�ҩ�.� �1H�]f ��7ˮR7;ľ�t�B�I<��3Uq���⸙{�S����WoA����X辖�&"rJ���!쿩=*y�f���,P�����y5�8:1�ܿg�r6
����Џ�e�I��B}b�om�� �Q��˃�z��xWe�aQa�AY|�$�3�`����y�h��������S2�����:x�^10��i�a���e�z���v�O���@5�8��dg��x[���� �N�,Q�U�bqS�j���?�*oR�Gƛ���ס�ggӀY��u��<��w^֎g1�L��2�g悍]?���2�?�nzN(�*��A�TM�V���M�Q�?qS��[8"α����u����ō-Z�6���f&����@F.��ڋ�Dî��Ԫ��˱��~6���=ʙj9+�%�v"NJ�՛� ��w�T��@I���Q3��2��(�����h{�nK��C��,��a�G��F�W�Z`rH�Vz��K� �cZ�'��*��N��H`�R:�r�<^h@���f�Ϥ4�Ǳe��h��-uqSS=�'^�-��SЭ�֌@;G��?T���HR5iS���ـ[��~g5��&8�#C�_�O��������C�b�Մ)j�"���e��N��}�ϝ�"�zl�w�=����l����HSscIX��]��|k�x�]��ӻ�)ܥ����]y��RS��:E��+�Ɏ������cei�^�c�];Mt��R�)�����%y��4�K��y$�~��0b��5��2޻`�I&�����&:Ć�!!"��6�B�;A�ВGߦ��hr��=��t�]�[�]� 1x�V��ʧ�8���7�������9�U8k�r0�X��>|�yfZS�k"��a(>Wo�`��j�zmX�������r��/���� ]yb�Ã�n���3�����/a��IPo7�w��T�WV���}K%O#��O5�W�s�nc�`I��S�m(i�E�e�A�k�H6��������G¢��q�y:���]����V��7��[&6����3�x���S'���p����'��p�P��F y���̋~���-o͔��N��~�WYnd
���`���I|4#�EA������qmE"������a�$��PO���Yۏ +M�Ǡ�M�!PS���a9�Ѕ-�� n���r_�W�f�#'Vc|z�y-�T`�m��ڍ!�im)��������Z�0]Z�Ȯ����8�������K�� �:K'(kCa��,�q���%ߔ1�o�
�����yg���=����2(i��K/�W���2������VʥQ�_��t�6�2����3�M��][	Xa���X���*S�h���k`z.݆��y0zL��u��/�6\p/�����"�0V�Y�Zy-�k�Q�+g���@<�@L-@���͍R��jU�����9/&���GC��]��<�;�
��+�JY��oM6놆'S�4�?�`�����O�����B!��7���cm2ud�pEkJl�(�T����:h���aq~u��7ŕ��q9�PL*w���;ުJ�C�{��n�X�2�J��F��	� v�_���O��8��t�
U��5��p� �7����y�C|�:�\�4 2GoM�Ȟw�Hw�����x���FF-�G^dq����m2� GH7�򵤔��l��@��*�I\�3�N�
w%���c5��,��j�8����I�GK	�;?�ć]��/�lTW�S�?���Cגk!^�~~\t�(�&�G����O]-?�������Y�5����N�.b�b�g�d �fH�l������[�l�A��*�����)-�|��7�2�S�{��a;�S�P�������1�*<~�����0�:�l�¥�12���6�@>���p��Iwf��,�$���B 3��T���nHE���iZ��#	V�f���@o�S��'#1�p���5���fԣy[�B���ɳ��ҩ7�e;��f�l�{Ve�]W�yr��p�蒭��{�|��S;�Y'�yj�9�q���_���6�+�k!����Ȝ`���%���خ��<�Deek�r��P@�a�&k���-Ϧ��bHr����G��@XA�kS��ǒ�;��
��j�W7&�#_ϒb|���[��d�ZK�rr�<�I��|i���Q���@�Ό]%�$"l��e52��L�Ȫ���y�M��&<?i�?���fF�D0OCxAډZ8�%�K�ʆo��S���N*Ppg$`�
��!�~=Z��%?�2�˵V�������v�j����$W(e��魜�#nBg�J��]H{M��/�@��>�X�b{� �`���G�D6�lbf�v����Tҡ����ux�u���jb-�w{��I
�v�*���H���c�0#ah����1?z��5������ry�n�]�N)�ckta�>9��X�Nc��*���|������K6��27c2�]���F8���X�����2���fŏ��p[2�0�д���&{�܅2��2t���":(���@z�)ju�G��Ȗ��X۪_떓s���"�bJ%/Wί�Sc%|
]|���U�>��z=~"H��M�ԥ��iH�/�"�ŝ�Ct
P�3 ���_f	�_��K�����;09+IZJߵg��HH�ga���e8zVV�%L�q��pQ��aQ!���*��5f3i��tvY-�2���s�.Ѻ�8x3���K�7��y����u�Nݽ�������D�%�-U��	��O��M�3tL�1iVf�Z��(������E?8᱀̬�xNǱv�����/Lt��.iq���ƨ����dmYc��Z���A��ِ��=͖��Â�'A/4h�H��_[Ŭll��9���u�ACJuO�Ԅ?s����:�r&�U�7�Ĥq����Y�S�.{�j��6Tz��T��T�������	�m@�U&lL����3�6&�T�ћ�]���b����Zr��Q��]+pX��"C��e���/�}w���2s�I��*�|�~�n�Y�̍}	�*��D��r�9��E����ʋ_�_�W��>�(��/���ж3+�J{�{> '#vͽ�j����$jm�5
唀"5���s�ϑSa	��+Q�㺮8Ȃ�� �ګFA�M�����虇U�
D4�ndWTff�$��n�r��6m�R'�%�d��pxF5����G��y�jG�0XhE��ZY?ݞ�Ň�O�Rx����	!�T��AE
��?�ZC����jȧ8�0 ����D����F�+K�Õaݕ*[4�z}���x����;�`�aY�Vm�d)�/�b;t�A���G��z��]�SV/�����BL�MHxӁ�]�X����M�BÔ�Mq�h��Zr6�������#j�d➡8aN*�z6ܶ[/T�<��BW�x�\��s�����m�ɝ�ӃdA�����w��o2�~FC���)MEzPB3:�m����IO"��@��U�������|o3����!�~吶^K7�Q
������;a�/�[�N�g�����F�����F�(��˦[c�o�|�kHK��z��9ʰW��?����I�^P3��
�)`�=��\��<��諎�c����P���n2Lj�/��K�-��- �ܓ}q#q<����r�+K�������͌:�F�T �_S�A��Y�8���+�P�>Y}�g>Ң���!\)�>�l����G��U��&paEI���� {��QNU`��]Y"F�<R��g㹠��t�M�fp���
W-9q)3�/_&�׀�`>l���d��c�:�j�Y
�:����dz'�N��B�ϥ�rB��4�b����_��xҏ!��F�4節ն��Bw�5Ȝ��M^f�8�C�0�õ9�(��@X��M֠�/�K/j�*���]6]�G<�/�e~���<����,�`Y�ӵ6 �g}�,�{<�	��=?�ɽ�!�6eSx�.53@ ����P���-F�L綊����j:���<X��u�M�	�r^�4��1��r��B4Q�*�����gǁ�-ǾW���.&/�}Ę�T���vEb U�z	��^vߠ�F�t��iX�e�#Xj]w�˳�t%�!�(�	,ɮ'���2؃
&��)j��9�l�!h�O��h�h��L�	�\4�o}CtDCR0?��=��Gr=�b2j��cW9�����	��˖/����������k��� ��� �o���R�����x�T����t�AbH4��b��8���%�|��A����~�pY&��##ʼ����L����[
���G�U��Y�Q��'ی@���B��pv �
ы�a�@�j�	;j�0Uw��x�</�ZmZԴ��@Zzv�`�<�����K�c��a5��p��ۡ�ǘ|�
�\�I'|5�WL���A}���׹��Y��/9��|,A}b�0g��⒝�ۻm[�}���XQ7�2�����+�r�g#����H����rsa:ק��Q��
�e	rQL�n@
��E�!�W�/���4�B�}4�YM"�Y�����o�ac�X�j����:�Mf��L�/� ��J@�?��nC���W�%"Eh�Ta��1��I�e��2�w�)��rq�c�r���S�>.6v
�
��&z��U4�L�������	vo!\]�s���Pyb|Q�}�����>p=�|(ܻw�Њ�/��Eo+D¬<�{<�F���'��#�R�3�1M��.)FBT�jP��5�s�규�'�=RG6>��wo���J#�t؊�8dK�}4��8�V��e���m5�N7��C���^H1_���w���2����<�n�x��f���bT�B�X[ej�^������ž�1
�6+ ���Э��(�W���k1g�*�IR@�������&z�x�8%�C�߲z�s �Yޒ��y'`ym�X�.�e�����B�b���C��vݴY�į����U��b����B͎�fv�-�[��-T��>54� �����+���el �:������/�eZ��Z�COs�8�KFi?�Z�������9��kV�?��������S-�dB�5b�|ӎRm��B&���
E�|��OU�݊���[�K�QȰ�8�+��o�������f�_���;�9◳�>���X	�!�*�3
�S��;��hÖp"�/bȔ��bGVp�I�3��^�:�Ѣ��Z��(S�\`RXm塺6�u���=ęh+��Y��0�>�y˧��Ԟ\��յk�˲`�Z�[�4`˳��&���M>&��~ �G�U?��D��3�㏄�@��Hᤠ�Q���0ͣ۶��
���M`�̇��K�{cK	X5�A�+ߐ��J�\cr�j������Fv�N����Ί���;n�=
��ab9���`�ń�#��(���qHn�`�P]��i���N�d`rۧ�{�6�5.;��m���ք���l�-�PQE'o=,�>۾	v�B$��ķ�-�M�H���e���'�2���	������κO��^/d	Y��������
$��}V|))	�!L��t
��&�m�X��l�2�겤�H�]o�,��ּ|�m$c���n��i	���U��u��B�!�"��{Q�ҋ�*��2B�?F��|���Q>m���	R>����x!��G�&r)�k��C��{��p�3p�Xy��Z�<! �	�z����b�S�_3�A�v�+N�޽��Mu-�7$k!;փcyoU��qV=:���e��9����RLI��'Ut̠ ω��dT�� �&�ޱ~�?'�5kfv�Y�m�d�YEp;���c݌5��^=�F�ere]1���cx�5C���#e�e������OK�o̝�{ڜ�X<��Ǳ�*{������	���{���"\ú�g�8�q-�;}\�	��3��5 S��3���!KR<`���o��W�����|�5��T�" �%$[��qѫwjSy�,��s�;���<�UT��� !Q�"{Tr��G'�IF8Өr��������"�Qu� ܥ�~|��<R#7�1)�E����?&?sz�畅��@-_F��$��Y#̇d��豀� �t��'�����$]"�]��!��0_׏��1����˚��5�KG�ΟȽ�W{��Bm��2�q,֌H�i�vC=�&Q9���s�dx�����w�y�i����f�c�g�-/�eI3uu)���`q�Q(��9��1(�O|,^�{$��.�(,�����
3���d@��S�>6���o-�V��X������[Sr�<������ݡt�p�������5�����W�|X�Ν��������zGE�� }e�w�iM�9����6�Jo�ɔ���}v�G��L��-�ؼtME�ޑ�j��@�m(U��������		�`��s��O;��	}7����#��ΐv7�ְ��y��k��b���գ�x�ׇ��]"�6��(#*��_��C+THL8�	Iy�VN�k�Ea\�E��4���\��V6>�
�gy�"�xϲt?���I�n͝��c̩W�	��x7��S��#�����+��`�M�˞��gd����}�⬳���r%��0n�5�Ip��?�߮%� i��Q����� b����;w���J�}��%��
��ʒ���L(�oW��r���_��٘�OP�<ec�[w�\a<����:�� �XәT���;��>�p�-ԗ���'*P�E j�<l�  ^�����U�g9<j	��j����\�!pZ�kN���熆DTx��qǚa1[4���չ�hA5��T6����7���p����;f7qaUi<��ˏ��2���Q���To���E��ƀ<S!4C�i�P�����#oh��Q�O��>�R���!y �k43�wf�-�n	�+))�S�u1�Np�9T��Pܒ-HsS�m'�C��)��(�� `~��)sp�RH /А�be}���6�tRm)_�]�fc��b�=��B~
�C��Q���bOi�V��Ѩ���B*�M^��b+�̮@M�:���(o��z�!�sDk$/�����cz�!���7J����J>��%��v���*�'��ae���FqƧ8m4'͸��l�O���h#��ؒ�����[x;2��h���/�a��cb��%�a�~4��\e$�'�Y�Ӹ���:V#��у�.�D/;s�.��6@zcr�*ܱRQ@L�'��!��K������I�:R�L�m���<����Fp�e\u`��?�p�
���	�ڤn����pJ���H9I�tn�
w=�KT�.�m����Wq����,�M8C��b����ѭ{[
�io�{m��0 &�R
 r�ee�T�Q����u�U�.�(���?o�[[F �(5Y��B�m30#�`@�E+)�	�����N�% ��{��dKd��\��a8�/�*��Ɠgť\\�Н�w�K+����Po����8h�����N���`4��Y��k�@��\Qț1\?a��=fk������W��d��8�^�H�@t�`e�2���a����vas�٠3i�l�܌�W�x!,����v�/��|~�-�����E�Ə�]�;�O1��B��_Q,6̭��f�.�б���p+�Y �v�G�m	��a
I�,sD�����)�I"���NH��U�](-h���#�wE�.p�Sį �n�(@ݽtP-��j�PBY\$%.*�6!���U���Z�! ��8��|h�3��M1VE�)�4��be�ğ8�V��p���6C^�c�Ş���3���|F`��/K�
�ʚ�������R8tZ������p�H�uK�$5e�.ٖʯ��.��]��2�� �l�<�%�\�09���"�Q�����M@��T��HZ�#1�X�!`&%��=�p�΢�C/o��z�(x�*�3�����ˤ7&(n^P���짞�M�(!��[���yc�[V4*OA� ��X���9<�'�,����F�N��T7q�%��Ye(�.��9�a��Z-�������Ɛ�S��*�2���;�!a�e/ڣ�oqz��JQֱ#�#]�e��#E[��4��d����^R�v~j��#.��%H�jΕy��e�Wq�Q]��N�w^��×�
��8���Tߣ�>L9��� Q�
�9Ջdc��2̈́㥍o��jY2�\����7|�+7-�Z��`��+��%H��"\=���ӓ�E1���	��w�c����koE��n~h�R�3�s����+&P��� !������{�̶�`D�c����+V�;i�@<&
�0�`�/�݊�Ό3���μ0�!	~��� �"�R<
�y˫���ɞ���	�4h�YSΒO���
�����j��/U8�2����t��[S��j�:�0ݟ��~�yj*�@lVY�m.9���w��*�lc��� 6�NC"�+��-�ns�It_'r���6-�[+Q�W��rQ����i��o(�"�w���¾ڷ����G?@p����R	���l  �(��7~�;!�e�;As���z%}dtQ�=h� �4(D�QK��X�h%����X�h�mg���0�95�$�O^:XK
�]3�����>ⓎN�>Z1'޿���>E#����`��ޜ�R�w���8��G����v���`s�,�����0��?`.3*��$Q�:�T;�o$��Β`�??�7��,88��S�r&-��u��ۍ�ޙ]�$�0Bb���{+z�F�c �{��//�~).,�dky���ᣠc� P����Y�ś6,A3(�����Er��5�ذ�{�ғ�9�h���CW����m�����Q��:��b�]~,SntGp���؄��������#φ����!cu!����/�� �i���?'͵�O��V����ͤ��&0Ŷ���Q�
̱_;��F�V�T��d��9�A�J��L];[(�ZMG�A� �I�r�<-���UM_��i��8��㎛�v���v�'���x�Z�hhy���yE� ��d׷�_H�鷹�6#�g�NTI�$��}�<S�=U���ո `a�\d+8T���^�t�Nn��Q9��v?�j���IG�ȎQӌ*O��o=Y@�����g��`���o�|)���U�6m����a���2�^��9�{�Dҵ���.�xN/:�n\D�Y&��eWh������ ^��1��+�R�Җ"{�� �����U걵ʢ<*�'�2Bmi���U���҂?���ɭQ�n��	�:��bo��TG�I,�y�=�2.)I�/�~_�4�w��_;���8C��M8��Z]Y<��'�ŒX���^m�Gz��M[��Cn���x.�z�s�۳����.�r�[�,I�h�	�v�Kd��f������X�1�����_�5�q�-C��P�E8��ѭ4��i�(�\9�Y��xl!�N��7���ӱiړ�˓�����C��3�إ�[�0��1��#�v
1u]�~+D���/��/�䇙�巔�̣Ww�K'�k��1�`��b�1P���3th�o�r>3	|.X���q�i��E}�d�5�reC���H�-T�p��[Wp�>�����ڵ� ��q�����6�����fUdbdA1�wThy��f*T6���_i<:%)W!�.�����OaN�R�(D�^�}�\Z�}5BA�ny'���Щx�6����!0C���[ƍ%N�ت�D�2������K.��� f�	�V�;��Sr��Y��'����k�S~�����˴M:sv�zHƧꄐ��mح?O�O�IHA�����i���K%Ӊb�#T�34K�P��D�k�N�)����v��xvH��P�7YO�w&�t��@
aH�z����#U�eO!j}�M�T�zQ����y���(=���l��������,�Ŧg�����%(19C:�B�PSxzy�1���Z��/�4�+$N��X�n'X����a�P:��%a��tB�,M���O]��;�B*��+�5z�>�`�����e_U�B����hʤ��B�zA�M��e&}'	zr��Had�����P{������Ã�N?��O)��Q0EJTV}'1���y��~f-��ȓ|IO
�O���3zCa>_��8�K�������v�vtl���y�N�u��lB�ｉݥ?I��j����!�,P�Kp��ʅ�/_-=��ZR1��c�l�Lp��d.\�
����e7�i��hX�QG�t���޿�.�xo֣�e�YB=�҇�gdk-eVJ%��F�B�7���V�7�a�WaS�a9���ˊŗ�N^�8�G��F��x���^����Ȯ����\��uF�^�	r�0�������?�}l\��$C-��"i=�鉓�� ��N/}&^_�k�ғuZ&{W�NsY���@�`�H���f������B$�W�����Vu(���$�t��y6��H�Lڍ���>���ݐ�b�]65�\9�*�ﱄ~����T���P�ޗ�(2������w�Z�W���#�*�̶OfgG�Ɂ��Ҹbm���͜T�dl�Q���H�3�(�Ψ}���t߬�Y�^��)'��@�@K3#*O�m'$p�@!�y��=
i��8I;i��b�}��~�>����U�4<¸$ЋYI\*Q? i�E+2@p\^З�j��Q��n���F��$''��v%�^���y�u��M,���ן�Ut2��&��0	#�"J����zu�19Tʙ�4s��"zp��j��YB�u���#hj'��ܐ��qd AT����1���̚3K��N؞�FE@���[�k�"��
�T��Bvo����w�Hn��
E;Sk�^U���L�o�'��T�=,��(��������󋝩[�󂒭�y���E��?�&�<��vv�+ͦF"Sj�[�
48 s��|�pH��Ô� v�t��೦��7�ƥ�7�0��D�&8���{��[��8�<��M��CB�@Q7�؄,>7~���0Y�%�9Z��4�
ZAv��q�-|6
���+��7x�Z{�P
z�H�ߕ�ϣ��(Dy1i&qn�-jN�{`���1-%�ܶ�l%��1F9��MW(�3u�S��+f�V�m�xA�4��}c�҄��6E��� (R���Hh�!�V��J�y��\<Re�y�'ˡC:�����s���* Z>:1���k����C�q#��E 54�~ ~��!D���q !�2$H�u�s�}.���B��lq4�<f�x�X���g���e� \�Z��oO*���ݴ���V�xԢ#�����.e��kS�þ��� 奴phg�l?G�#�6���Z�p�K�G�5l��?"X���⫷����e�/�vALt@8>�p����OU�B%�o��D�ߓ��dJ�_'J#:c+ٚ��b���!N�����G,����Uc�%�dcC��-�Q�E1���v����hl�>���-U�"g���1��O<��P��ᝡ��x`Qo7�)�֧�X�~��>��{��ܖ�h��a�V��&��f{e�v"'G �XP�sH���Xfuɲ�x�B2Όxeg��YWq�zi�+TUy�w��tg��ATC�}�"N�)i���G4��Y��q�M �h�0l�( ��ν����ʑ�"c<j���gQ5���]}g*$�H8��0�3����k�V�ͪeN�p�?{�@�U���͟����i�����Q��g0"a��]�\�>z�b��x��'��'<��j/a��e��X/H����X�X����K#���z�&w�����{�*�V8��Ll,%�_{�*�*�7���q{�Ʌ��Z{�[|��fc�C�ӈ��NʠEʙ�z4x��q��Re2H��'�����@>lc�-5C�c�|�p�~8��Xw��<z�����c>�3�}j��Rm�*Kw��X����Y3�i���%�7s
�,'��f�U4"�������>��
W��3~'��R������уx�q��o�����C�ڼ�@W���o�e�FX�3�<b��K'<U��꤃�/?�� ���
UN���w�+M{�֫r��=��n��;5��6����}C��(�5�DX���t`C�o�^g�L����4��ˆ�]k����Ǒ7K�*a����C���;O���Z{O����㰰��8G�ȷw��sL5=�v�(L�U���"i"(�}"�Ӂ��X_:�+!���=~���k�u/�7�gl���j���h@<� �K0��p�3c	���Gl�c��,ҳhG_�y�v04L�$D�ߚ�5\��,������؅���٪���f���j�S�{�2��|��W��'�T�;#L�J��������]7�%K.,JR�KP�.Q��Pn��۝yf���jː�Ӑ�7����e��D��*��v�>o�G~`[`�����Gi׀���v$��bm�,<��6b�[�S�Q2�	ɭ�YZ?�L Wh��%b��p]Sa�����
� �զא��Ё$��TB�ƻo�uK}��!af v-��!쓏(��D6*��q��Q\?�>��k�AR��"!��O���e盎y���>Y�?S�~���eK��-pwT� K��ޢ
��Q
v��Ѯ�|�ZT�2���r������*/��z�ͳ�Yhr����5��Ƴf��$�p��ˣY�e�ҁ�qR�Za����G���!�����I-�AC�g���
2����k�Z��@���E�':��5�I�|=���
�D�H�����ѮF/g�cJ),�J��;�)։j�FC�4'�K�h��|}�qv�;�X��ųp��R�!p�}:���wS�Z�!iI�3k�����|h��c�%t&) ��9�n*J,��'S�$?��^E�^��st�n��Z�n�WQavD�Z�}���[�(���9�00�pF1
X�cO`�N)r@��ʲ9tn���O���G�����R<�jH�;FD���/�ͩ��Ұ��Lt�������,��I�S#s���d' <�����JD�̇j<�-��/٦B�Lr:�J��wX��F����x�S~���6��m�IF�4�D
pq�n�l�Z�Jӭ30?C~+^�b	����+_cy�^@�&h�Q��X˭�5W�-N8's�F��M������v�G>�y���K�(��w��FW�B��-�O�
�=�K����VG���C���jsfk�@b�L��b)9P�7-����/b"Q�dy<ûL��� F��bto�jW���<�XOB���9FP�0�)t4	+��ҖP�s4z�V(`���캇������M��L��9�K�j���niI���#g�#�n+��X�� {�q�T�.�W�F�2.��Z��
m/u�V�ѽ�$^��k�y ~��/+i�oUN8��&B���0�[���C��j[ �V�z����ċ�:�SJBW�������u�RC�
��u�b0I ��3���>���1	4-ǘW�V=&���ږ�C�+)�D�6�Yaj�j}� Ũpٻ,�Ď�����IU�׮����|<����NR�b�9c������d���y*���ڏ2�o��Y�<C���,��� ۀҮ_4Hn���@ę����n-mv@ܗ�*G}"����f)V$]�:&��=
ˁ������E�<@c89'thJH�����D�<��q��Φ[J�n5�xѵ�[�m'7�-��P� �E��2�|NtT�{}|5�΅��m��D��4���lt��n����j�2ֻ�{�&�-�T�w<ץS�}�] y�<��yx�^�׎��G�O`�I.�����d�&Fu0���#}@65�1�m����ꊎ�b�O�Ca�~YG}GO�*1���N!��μy�k��j;�8yY̊��� ��~s$iT������vW,=��[,�K�K*��HQ$t�ї��M	���fԧ������PF�$��\�������?[�z��!\}��$N���n}&S���\_�LL�[�1jw_�x���#��:T�{Ln�=�jy�h��ir�w/t�����J�BP�����
�[�^��\RY뻶�V�wrd�^i���d��	��H:/E����	��s���uA#mc��A�K�/ct�'����DS�����t�S�M�xU �͜�N6$���3�WEl��)��򳌰�I8_hV�x�SMK	)��>A�S�w�$>��t�/h�5K�e˅W_�jRw�Z4�4L�5�������{,���Mrv8�,�s,!^�b|����Q'k@��:����-��P	������������
'[�2�x�m�>��o�炒N���y��Us�|.�Z�?�����B^L�.~�P���`a%�.�����p2o�ċ���T�d�3���PDz	.c��bS�L3��!,D�h��v���W{J^[�()�^�SX���Dk�l�A�Q����,Jo�ۈJ��]ʯ�O�,Փ�$'.���_��4�ʑ��d�N'�F�[��S�>�v��LW=���B����r**�O�ڻ�]��l�iZ��� 3c|�Ѽ`+٪2�����\�B�{P�D�S��k�I��c�Y ���R�P�34�ZO˭d&��On<E�	���\��7��{m319�B�Q#+8nZZlbm`-W�ߴ��~�ZR�^]���S������M'�ؒ�B^ec��=�������-���:E�7��s��O�YK��#��Y��3H��{��Qք��"�����TO���
��d��V��R�mBZ��d�1�B��t�p�dm��j�G\�.�>{�(`ـ0Ǯ��x��<m��.�|�:���I5F�hE�-��F��f@0it�x)	��c�Be/��cd�R�yv��^-U3H;b1��!��-�l�����ٓAC��>���q�@_F��T��=D$I���{T��G@�=�ջ6�B8A����7��l�JiB�-%�����7x�oe���.v��;��U�d@mrN��i�Q�1�?^�G|!0�NlS?Z{��{���	��F�gp "_;�qo��a0��9uKe��xܼ259gnw���Y�D��&_t[�3�v|�$%��/^�3�^�)��Ι��z��ܯ9N��5"�a���)7OX^n;�E��
���?�&\;ȸuױ���S�W��(�a�S��X�o>#���SRօn",���4Qx�UV�\x(�l5��V*���'UP�H�j�Vn`ɀ��4�Ҵ��R�M�9Eh7�ZjΠظ�R}��Wu��M^�3㰁�f��5HA^q�ɾ���e.���)�q�N���qvʞ�}�m�Yh�y���b�V�|T�i8 ƻ(5ɚ��\�L�uqm�>�j��������+	�N�+�my=Z�6o�5�%��:2�f���~�!���@O��,�)0#5�iP݅jQk�畍S1�Z�
������W>p�(b��[cS��!�0����w�������24?�(ΟG��Q��.�Vc@ǻa`�N
��F���%��6k(�HUC@*��:MQ*����U��Hp�/72Z�k�u:ͨ��"��'�ȿ>>+�MYj"�>a�A�������O�k!ê{�����ӧ�C�?�cնjV�)z�35?�����R���\Gm��Y3�dUc��-�pP�c7H��.GL��4���
�;�>T����|z��<�碁�S��)���A��4]V>o�vTX�	)]�����T&�蕖��� ��y;y�:����Ic\����ܢv$��E��bL{m�m!�F�-f=�,���Lx�ܚ�O�ԕ����;BL_چk����rR)����? �;��mi��� A�J���~IHR0_��e����)�fӂ9*����( �m��U@ T�Ԉ����2Hc����7�"�������,eJ/�p�m�#��6���ܽ�b	������l6�@�l\:Ek�-k�{� �k8/Ό�M�[Y��W��k��:1�앎_D� �_���i��YA̓�	�*3�D�r_$Ԃ�Ӟ��]SH���n`B�1� �D#�ws��v*e�r'�p�6iO�� +�4]���uD.U�O[FZ��?7\{_�J~��]3��~sD����*i���j�i�l��.��X��Xӗ�\3�-1^A$��ť�僿����^��љN�x-3 ����"�ƙo�ʖ`u��X�{xZp�Gp��j˖r�tL�`Iw�3�`�,<��vQ��`�[���v�����D��r�y�:�q�T�㇣.�'����XӤc��{.�Ed�͟�Q1!��Im��V�_.��vkę� I{n�ʟl�xDm��+�&�{?E���`j��fu��SƊ�F����t&�P���e����Sh����2+�Dn|س�Ճ�<�EM�)��r]�E�E�T��@���f�շ��e�J��Ő�(��@B覕x�_��E=��&GL����"���n��Ѻ�Ap]�u
�g
��f��:�"�E�>hNb?#c��P̠�>���+�^�@B��%���~|h�[�%�ٶ��,U��Y��	����U&���mD2��\o�M>�WR�&�@|��#���ɿn ��Jr�9�����Dc $6EjqцW�it�ue�׿D�SSj~!��c����қm��v6Oj���ُ]A��$Z��@����0c�����'��b��6�M ���Ìl�d�Ȇ;4�^���Q�ǳ3.:SlsX�(�60v�Y���L�b\&)K/7��G
�h^����$�p�����k���j�͡P��qJe� ����+�0͜6�궚�'s��+�Y�B�Qy��!$��Uz� ��Ɩع�!:��s0uS'�ڻ��a,���K&%���-���II �<�_�2� T2z߸��瀩�?9���J�@���뗔v��P�J`��I�Π�W;�}���Ն4{C�	Yf��MH��Q=��E@��װ��g��o�(�xgam�Q�ύM7k�=ʴ���G��S��Qt0�)�)C?�	q��D�@3�Ȁ���E�D�<�������X`�d�^�����{������<�8k���0乫/Ѹ�U-��pnQ>�2j\�h� ,�u�{îܹ�Mл�x^;�T���+ ��oEBؓ��9��^Ze.7�8&���/w:���8�ңiM�!��}rz� �E{��a��PV�W����_ai
H�����������!0~�uSl��F�z!��d�
�Rۺ���K`���'��Tp�5rH����i�ƣn"z�\��q&"v��hs6{����T>O�	G)#�~E���z��e�.��=rG)͹���T�����.6��L_�������ޖ|v�0�$[)Du-��isC�C^e�,\�Ѝ9o)w
��m�J��?΄8l>��@��s�zthO����|.�b̓k�W؛4#�)���?I��2�a�5z�)4@f��~_`?��y.�V�6)>�7�.�_�7u��P�%t���FsZ�r�yNIy����T�p�8�	�t~�� ���Wۍ97l-oB0(?1�!\{�\�E�0g%e����
��_9hv���;��=sˎ�j_F�ÈM e�Nws>6\��@���B�	;c�禎ko�����`��A�6Y�!z���g��>�b]�C�闿��Ħ��|���[��(�����z�RͫJ�����)~q��_���]U��"
�%�u��dɣ����]H��X��#:���n�H�F��>����� �G֓�e5h�t+�ɦ�=��}SKSH�B�mW��Q~�%�)���Yf<���Z��[Ͽ$-.�#ȫ��v�
J�͡�Wc5n w�_)�^�x�|����)��M���T��{��l�V7�W?�����pC����Q+�[/ը_�����_M �W�֗,�u
�462��������~�m|gXϼPx9���Rq����'g`�:0�[���ͺ4j�{J�-.���{B�b����c��ot�ǈ�B��wojZ9+:�;v�8���&�U�i:G#�c/���õC����,�2x�9;T��&BH�9RJ�(���?���q�Ujs�t��6&_�|$��и.���� ��ݶ�N]U3���$L�8�W�Bx�4p����{�i(U��|�K��I��*��̕�J��y�1���>��#��A�!M�� G8\�p��ΰS������L��t�(&b|d�w����G邺�6�Rd-Z0v��s�!�Iz�]�Ym#���
J;[���Vz���G�������1<���T�ol]�L]�l��4++�׃`r�6�x���$n�`�Ĥ�G���¸_� ���ce�{�f�)�U�MӰ�����B���l����P����&)�'ƝN���WSAcsof�؇�����=���=;=TT�*x�`�)S�r�-�R����P�t@���m繒���DdJ����]�0�]ԍ9.鑰�o�˚<���P���:^5�C�������3Z�����A�H {C�5��O���xӀ��F2(��Ń���j~5��-y_�Y��A��I�������+��"S���<��U`~����@V�~iȀGH�A�y�߷��
��b����6�E����l0 Z�Vp�V�>�PaP`��4�k�7A��|z&\4O��IG�{��,���<�>��(��E@�v��ĩ��� �8�.�i�Y�,�&a*�1�3�_�鱞{^� S�� ���1�҂���k�XO��`=]*�� ��h̞7�(t��C�ORP�$+�p���k�k���	�3���Է�_Hg[�K�8W��A{�r׈�<#��+���\���"?&�]�L��Ln%:���ZkF0�uN�E���Kc!cu�<uу�`u�U�#��_�ޘ����K3t(�C�/�m�\�N�����f��}����r<;�%��_��U����S
��[p[�_���>�0��Pg~~AT�98����I�M3Gv�JZ2�&�/ο�@w�G'��dm�=�6�p�t�x�{#�+dޔ��1nZ�^?k��mEd<�eR\F��8�M�yN��x�������ڷ�v��Җ�LKt9�n|��C���G�?�4����0qc*�X-�:��p'C���2��rD!�������uq�<��2��9C��`&j��|G�X�g�u�QID��&A���9�Up�+�yһ��g�C��]!�܍q1]03υ6^�P����f��6����-���<o]�-�����&{h{E���s�F��\rl�8�դH g�9H���z������'�^�P�[Q���@�� ~�6 �C��s���aJ(�>�40ø����r��BS�Il��&���=��<e��>F��\�JO\T�g���C����ݤ':*�m!�Z6�m\gۑ��DoA�e��}0�I��K������򾽁Pq�������[	������8� �^���
@�O���?��Hܖ3���k������.�6�
:���G���eB��B��Gk΁<Q�8��o38~�e��#�-m �y5O�հt�d�8�)��l���7�}�v��N5������D�>enꀋs/�r�-�$з��������?�!�H�L���;_�Ek'̹tW�ݭ	��Y���}��FCja���_H<Qkd7�l�����k��"�8֨I�np�b���z�z`��4.sp��*��8�2�(4���+s6�0ЉbGy�j���(:���c��E��j�3��?��eQ���OB��:��̗ikW�*U��(m�/A�g��> �O�Zz����4ٕ(�K�5����\��vsP"�c��m�Q�t矝��.��9V�O4Q8e�:S���dW�s���`u�nK���i�zC�tS�i��U2p4�B"H=��(,�cq�	�pgBk�<sր���1e<j
�ۂa��w�o���9��M\7�q���Ut�9"`h:~dJj��W9)N۲�c�;�w~�}�>,m��ی��q��� ��r��M��n��q��"5�(X�a��4�t�7�/�Q�<�	dPt%A�:k��}��#��J���i��q���`���̳�9�h%bX��;�DT֪��k~���>U�om�v/�ɻ�+K�|����h�}�UY!t�o�����2b���Q
[�Q�f|�1�](U�(��]%�������V$Y���݌*l�e�]�.C�R(Tw��hіK�{u�2G�)P������wȡ~��<��I\[�0�����k<,3��m��CZ���-����0��'B���6��ݜ���$%�\���� P����3��I�yR;�2B0ӟ���0A�_��+-ěω�*l������[ޏA���:��_��P�5���y==	k�@�nH-ؗ�Н��a�<���M�ɹs���X���ss�`�pyM=��8Z�:�ۉ
��e��o�'�X��+���B#�=���h&��DKU�\A�`��&V�/���nVy�XAƥ���Y6�~��|�y�n���k�#n^7P33L�����\q�K\�ueH���� w6�¬�:�["��H�$dtA�����z^�]�5�!�I�6�O��i?�$�(��v�ku�(�O�����ȡdy��FQs�.mRe��i�Cb�>�7�ŒX̩5���>{�0 �>p__��9v��
�'_}�0�?���4`3c*�1X�.�XG�'@���"N�}n��s�l�oh�ڜ乼��  ��ȳ�0��|C���s!`���/#h�Ƶ�w�@9�����=jɲob����4�^4��,Ih2#S�@8�l43�.�&��l�Y��ŝL�i�b";զ5�T���YPrʲ6����S����[���S��;������qw��J@��M�	n횟�+�-�4��Ӛ)���lg�  ��l��e������<ϿOa~R�f�U$�u'�h��,�2#���Z�T~uα99���q[��#�nb^A�A'`.|�u�ǞXi�u~����[C�h�٥��D}�zNG�v.c��6b��X��0GO!*���˨Sv]�ę�P��>�SR��25lju�w6׻���E��
�KO���d�ǧ7��;�}�bL�i��-)�潐�xS<�5'�RF�����(k%&�����D�l5�*q�L������s��˵8��J�����bb������V�$S�m�����&w
n���x������V����_��M��75����U��4G� �b�Lf�Q���Rg�
7h��~���4p5���F]`�Ж�jz:'�@��iK �<�J;�Ew0�A<1�:NK�����,��)[M��Xa%�/��D2po=�W&=ۨX]ϑ�ڀ߯�3��Y���/1��E��ܺ�������ᜍ�Lu(�-B��J�]<9|;�Љ�C]W�`.�p�~������d��G)��<X�n��a��_�	;7N�8;F�	P#�1��72�D�,n7y:�w��D��	*��u���J��V:��]��{ȅ�v�U���"1��v���&�~�?�-#逗�ゝVc6h@Ss����2�_����ʢC�`�X(�B#��Gʎ>��L��:ClԻ�D"l��� �(����8m+��W����&4��MLR�w<�՗M2�q�)^��xu��C��9�)0��.x��/9�۬���G�T��G�$Q�8�]�n���arɚ�ʝ>��N?4��q�D	ѱ������4+XT�����g����K�/-�NUV��Z�C{����Ҋ�F��Q޳R0vֽ���(��B5'�e����օz��Vy�C"�g�¹����5I��#�NWR�����5���4��T�!�QX|�^�g�WFRTB�P>��/2�0n���ol��0�,�o���ƥ��Q�0lwKL�^v5��4A�����Ofa�MJ󞟍�q�{56A��]?@<wn!�gΎ5��N�eUڎ;��7�I΁6l���+;�q�_9����jƳ^��'@ �&?�T��o�#��K��R
���m�9��*9�>:��x�t;j��Lg��k��3��`:����KGW�	*ΐ,�g���8��y��NM�C�cNn�k�P�k����{5 �7w�t��|J#X�Q�%���g`��n�G+;�s��X����M��?����;��k����|�f~�{q�^�Vh"���1���ǶR��v��E�RA���>Sv�r��H-!ץ�p.n�z3YV��G�|p-{�����\F3������(Y��2b��[,r�M��G^�؅���صB�i��V��V��X_�(1�,9��y�t}rAl�| N]4AT��������J�m�L�{�Tr�-��ͳfj�Ɍ�c��𲳍� c-��Z�	��?�4��wg�d����&�$[F'�J�E�|bj�����i�u�2ѽ�}xHW]�P2��þٚJo��Ԇ�!�����`e���_#��He�'�����D����Ծ,^$R�M_��ѱ�gd�m���(��J�[�y�xW烢e����E��;��si.��|�D��S�*�F��I��@�5�5H��2���f��SVK�7���mﮒ����:s�yr&t�A5�e���?�ƚȷ]���P�V6.%R�J���iWWm�ь���h��s����/\lAރ�
�1�x���B���D�Й�v]|	V�^L#�� ��$t	¡<Uӄ�7BiwI8�pg�*���r�^z��10�܂���
߀t�Z�\O�}��r��D�$�\�Ш�E1�F�L�8��o#�����ZD�rO���#>�΅�$�k�Ϗr"���l���\�HƚX�!,L�jBa����or( Kʃ�M�.Wr�����0��_Z�hV�|~@��&��?�pI��kz �4*ܸ�ꭷ���c/�l��\6�]5Z̲��Rs��|���c�ȝq���+���h��	�I-�*�G�.�=���q��e���E�a-�!�ւB��Q0Ŷ|b��ʌ�,�q�\|Ɵj廓�d`X���:r�z�~	4�}��/~�.^������9��n��stY$vS��[j����Vd����8U�ܨ�4��^N�N����,
��u�R`���28D!İgzD�f�����x ��t�s��E5Ӣk�A>YE���kp�SǬ�@k�hE�P5`�˕g7��"ȹ����Q)ۡ�fq�,�����MjqCR��PKW�䴬�����Cg�F���~}�ƚ��I��8o9����[^��l�Lw����z$�U:Ĳ��?�h�o*��1y�H��#�Z����V�c�Zxj2�ȶ����Z��;[���M��W�U���ɭ�yx\ܓ�ۀ��B$�[�f�#q����?pJ}�K�qqYίAζ=��v�K�8-�U�1�ہ�����d�:>�x{�Z����M5N�	�o��|<�.�$�?k���?&��K&<����i�pb��ڭm�
��.�/\q�,�@�x� �Vh/�w��b��o]�A"F��i�����皎:����qz���<���2�K�6�@� �x0��I#�6���!�~a%]��j���bɻ��q��ؑN^�� Q��L'�K�gRT�`Ğ{b%�+��l�_9�Υ-���^��p��6{E��{k�L�?����9�G4��N<�<pZ@�hJ_�����W�]zn�T��T�/��~ȵ,ΈW5��vA�����H�M��r�;�Dw�xn��s��[����CCD����p�&�Z��T!�$t�щr���ű��IM;����[�7����$�S�����
�g��� eP4�|����cۧhH���
tD��X�V �oW��G�~��Ee���AP������EnD3�q�h$kN�dY�R4�=�D��9�$�/ʥ�o�֥#�|��ܙ�.�蠢/�=ro	�׈ӗl��EWú��n�h��������bO����@�F8I���$f,*��%��~��ͩ��$����D <��KK�aB�&6<�L��?���}�#vW����\��sc����~�n�Έ��K�<��Z
�|+���q�R#�愽�PF�{����P��t͢�i�ac�����B2B|�Z&��@$�$���r���ELmg�C�}�� W��D8����,v�q�P��}������q�iI�Eb]��no-��Ɵ�c�G�zh��6;z����Ȩ1,
�\
ȧ��K��Q�
?���5BO��J��:�-�LE<Q��؁��R�. ���P%)����D䝤�� ���> �		x�v4��}�<���=B��a���y��b�T�)��;�y�ÒoM��Hm%�<�S!W!���h�4�(n�U��-�w����N�u�P��CR���0���1��]$a�ny�_ڡGxs	�1`�㏇x�������Zǿt��U�\!І�ٟ�8�K�F�?�X��Xn`ϲ�gz���=��m�l(��̌�67\+�'8W�k��o�N/Mc����+�-�F�u7Bi0�h-V��Y l�"�i�Q~�2�U�u|:�t\5�1:h`h��Y��,|M%V�z�?���n��E,��Tg�ܞ)��p��F˘!y���d �
�T�x�t5ײ�����S�KA��c�rށ�ba�덴
���b����ѱ�a�QA��=7 �C��8+>�!m�ڱp������F����`[�k�:��g�*��s!�Ş��}d�����#A�!�;7J�T�IJ��6��L�Qj1�J����",���7��:#o��L�l�2�#�|�V���و�}֣ͩ�^�n�Q�@��:���P��%����r������r]B�9�����L5)�F�9�4Tk��\�^w&��G��]�d 芬)�k����
�2��HYl��[��~�z�[V��n:�f��CE<�vL���
�*U�4��F��儫]�Es� �d?)|�O��|�ĦN���a�T �#̰5�]B��⡢D؄o����B��o银ZD����P#��WC��6v���{��O�D�?�IS��(��u�Dvꔵ�#P2��:R�AN������&��4h��\�c�Ђ�^q�3�s�WW�x�g�96�a�'mВ�*_"���n�ЅG�(��x��8*��2c���Ch���G�y���SW�P���OW�qv�Z���q��_�g<��j�<5fBѠ�'rR�6b\�<IN+j6�f<L��W�cF����heX��p���T,rKx}}��=9��D�reM�=ro�3����I�/[�#�(� \�@��	q�x�>��.*f�aZz�+DF�SϷj�fR�wP5�-C\@]杪;G�J������A����
�r��re<�
l� ,��KDM��{��
y;:�����KN�=�� �Nb=�rO��s{"&'I��K��[��ƕ�҄������39�S{�н����n�{��Q�ǥ{[�;V����Y[��[~t\��0�N1R�G�yx�4�\RS�n�"&=� �Ud��Ы��B	�0�Ô�ɥ����&`�� �3�V05�������=5m�Jy�	��s�Ms[��$�� �r�ȥ�Lz?������M��%�W>�)QJ
p��矿D��=��]뚃\�w{ʬ��`s����S������͈�a�rY��5����,Q��Q��v�M��f��&���wH�a0�|��1��@]h�A���e�:B�AR��g�M5�u�k��Ǖ!�{���7	T����7k�{�7?* 4��S���="�Cѳ�om4�f@����&H}
 :�0C�����&���C�S��I0%KFzf5�m��?"R����3�J�UZ����/O�/f�;/[����JJA6"�p�LB����-�m�'�=Ϭ�
���c,������}�f���=�8ۄW2����Gur��ֈ�&�J�6��m��@� �`���l����[,��=�"t��V"}�&��^���XO�i���Y��Kş�V~9&�8b��Ɗ���@�{�/�{�લ<p���o����j�.ۅ���M>	�>�"�_Ə�4E�\��;Xܩ��.�Μ����������Rζ5�|�g�=*R'�8�\=�C�S<�~c�3C���`}2=�J%nV \ƶ�[��	��\�ɍ���T\A�t�� ��	0��ϾY�S	"*z��H�舉m�,q�2�FB�E''�k
�2���|��twZ�	��Q;�2�����;����v�,!�
��5ky+�r��c��y����"���&�Ș��`v��D��`�6���/Q���0 �O� ��b���z�,NܲR{7��l�c.[:��!�khD] (H�H�fFǓ�W�4ʒ����'k̸�K݇��vW�:� R�h��b����?�L�����v���J���T�\�9~ڋV�=l0��@#���������0X҄^j�o5/�|���0��<�?E�8BRY����� �[8�F}�{�D�l<T�+xZA6,b��>5���J��ܰӽ�sV=fK���I>���)c��S�A��X7J���z����L�B3�ͬ�/�Ȗ�Yau�=��,�'ʳђv��h
#l��U+r�/�K���*����ê���V����M�ʤȟ�����7��]]��ݱɜR枿��#Y��N����Y��j]��-�yz?�?|(Gֻr]��@!Y�]A=��4^[������z��p���.c�J-���u)36v��b;��dcj��7�q�R�Gܐ$�z�����;���e/b`����;�p^ ��j	�vEv�?�q�S|i�5r!���s����sHG�e�ʎ�Im�6�%@mg�>r�D��#���]^�3�/J�K�������\�W�ȀE~���QF�e�7����/�7��܎8R��˿�c���r!�!]:A�{DS�<���q�)�뼅{�b�q�P<�3�@3�_���n�Up���p�s{��R�x�/�『T�z���(K���?\#{�kV��*7|��^.m���&��\*1¼6��nz��[MG��)�Pd1�VE6m����s���<T�A?y�Kz� ��l\1�|t#D{v�N:;��"F����x@�ڋ#ʩ5R�2���e]�e��k5���S�cޠr�?7I��R�K�b&-����H��.���' �V�c:� .��l��z���{�����k��Z(��O�sN5YJ}�{;+$�f�����^kiw��T�=�c��B���@�ABm�Ԝ~�$�gp��S�	����g	���^�c�%���H�t6�#�e���Z]��-�^�'�F�x���$�Z�̔d�!�S+@�:��x��eLMb�^aǻ3C!}�;��r&�ze���ZJ��B�TCDa���O�d	�~�����=6�*�Z�\����(��恸��㐚x�U�E~�Ӯ��]t���Ek���R4/���
�/���^�^�ٖ�L�É牣�Z�����w��C#"����ʉ���\oq4�=p�\��=E@K�6vt0>m�x�SxK�L�,�h�� 0���3<%��եU���!&|R�A�,����X��vtͺ��j����5�|�1�����&��.S��\r��[L�s�'zA�(Dm��&�xS�w �r�7M���F]�Yg ���H�:�/���9( �/�ƫ��M�qb� t�#�$��Ew�����`uԂ�3�����?sI��_&<,��f��FU��.Y�(�jOCΌc^L��U�W.�-�ŋ�$���i���C'{�V�36]~�P�Ap9Y.N�
<l��-c�4�f��� �D7N�vX�s|l+A� ��Bs�O�>��ǤZm�O�� 9�0�b�P-��+���\��z�Qs���"R����A珂=���9���y�D��Q4�'��	u� 0�f��� �ɩW�@��0�^���5��(`ΞI���C��D�|E�uՎE�[����W>��6|��ɪ]�2�6Y��=u��6˝j*vS���>S� ���}c��U��$��T,LP|FN;�14�,Q��KtD�[��0� QB~�(���Z�yV􅳴%�0[Ըn�FBu^M4di��ԑ�}��s�W�^�����5�Y��A0LҔb���l�Mxæ�=[i7�L��i��|T�L�]�xA�O�]{����)�ڈCKN(H�	��>P�c�	*[�O������1׊X�������?���q%X@E���/eJS��q��V�ޡ�!'� �X��ߺ�|��@������,�9[F�]�������&bLҚb�)_'tn=��|���mőG?��i�W�o��ǽP��ܿց�O�F�T`7��B��rV�~��T[E�[��0	�pxt3���z����o�>Q����I&0����e߆O�|�B2�����s9,�yN?@=�
�V�~w�n���lk��%�K�~�.'����9W�?Yci�1If'����$��~a���k�~�Ovx�_�W"��M�q\B&�ᷘ �w=OP(�p=��f��
+�9Ի`t����U�fN-ׇ�&b����i�S������ގ1� �����;ܰ�w�R���v�e���
�g%���3{{�Aj�"�w��.v����68Q�L�M���a��H[�Q�֥J!�Uy~.���af8�E�{wv9jN4G.4t�uKP��W�*.PFqM��AlF���<z���jAM��O���	G��A��Bi�4�(���	^JabvrcDT�5�*o+����|��N�o�Q�3)�������f*qH?�q��Hb׳��,�}�[*���$���ِg��V��_����O�$�Ҟ��n�n{��v#tdn�;���┃D��>Ӝ�� }�.�����c&C���[��*4�<�jd�D�QY=y�6X��R/���lD���_ 
��Y��PE���џcD7+:��u<�Ä��E�N�7`�Fy�_��y�����������M�8��`�aWPqZ_������dc�/�#Ǆߓ�q(t(�4R��C��6Ke��{Tw=����x6��j�7�,����e3�J��e��5����������[0�U'S@dC�́iP؈(lU�<e�3A�e�m�z����3ϼw���i!��'������0h�%ݍ}_�}bd�NHX��Ep|]1��a3�c�W/c�F��C�>0�:ֽ��>��W��&��B�-��	[�:���"��%�J.t�M��D�:PE �H��w��K�$xv7,��؞x���e()�z���t�0�$\O|t����.�<ϭ����;��I���0�Vp��6�T��LQ��(����;$��A@�M���NZ��H�\"�",�"A�I��e��7y/~$�{���"��Cw�^Qp !�!��{3�9x�\��"� xv���P�춠�h�w;��@Cר�OP{�@�U�߅�xl�V�0�*���_��S���s0�F�-��a�Q@�5a�P����E��o����0[����QPh*�I��A���"��^/Yv�'��*yL��`�0=��ㄊ�]E���f��{w�]a �,Y�D��*$��C1){�[f����ii�wo����r	�a*"�;��>g��$�N��dzw�-E���d�ۧ����ln��p�� i��n���(.Y�2̣]S�	�1�sq"���j�`n�GA��0;�
�_<�B=�U��T#ɰ��`i�{�m�^ǕrŹ�į�w�p��ʚҙ��<�������o2E��UP!s���ԫ�3��w��`"��؆�Y��pZ���ŀu�����������w�a;q0��8SN���j�{Z���Cum�~bG	7�j#��9�h��!sDyEW�c"EV�TK�$��o��n�k�n�n|�=e�l��y'L�֫�a����J&�Ծpm��n�'�΁����?�jU;�� �KuF:�UT�Au�2��A�:y�5��F@;�¦S<,�N����b���Oė�d�5� ��rF%���KI�z]��h��2�R)�z#��5З�6��wuv��;���W�%>�����.s���N�8�L�������n�^|\�]��o�D��g$}ec�TO�\�B����לGC��0]HuZ��1@���I� ��5�L�»�W%*�F��*`�Ng�O�
B�Bۇ���Q����R�����f�*<� A��m�-U�_��� �"¡|�f��-J��ᾭW��`���:�N�-��D�]��X!�� A�>�Gb�6ȵǊ���C�ʹ|*[�q��CTrr�!�K/�r焆͈U��S�s3q�|��`c-A��w�G�ꤱ��7/ג�P:���/8�-?��!bL����5][Ԓ�} o��Ɨx��`�����
U����Z�C�ʩ�Ҳ��l�@!�������J���OGC���i�E�6Tg-];[r<l�c�n8�a����_E���$�"�[�~]���q��nO
ʘ#?�����>J/H�ߦ/�cl�Kw�O��IT@��[tr�F���$����+K�0�h���E�w2��^�R���v4э�Bgca����8]��鲊�	�����*C0ccP8�_(7��VZ ������;�Z�Z!d����3e��.��g���X0�;����)d&��g�ݢ�3��K�n������F���Z�ז��m���.��v N�a����@E��ccR��=�s]w���u���V��c�C�?e�gv�2e�C��t�"�,Ӡ�"�_�w>�|=�iȫ�'�ɝnN�/hf�&�G��Q�6�[|=��6ip�&EM�:��Pxjxl����@'`kz妉|ߖ�ϕ����GXvq��۴��B�*���q�W������>O�k�GB�?q\���~.ߕ�V���3k�L÷|���:6���S!ց��6�^	���8r�p��������BÀ�ɼ�Q��X����Dq�h��s���o�%����1��v����_��	|h}���=:I��kGc�%H5o&v+�
�CO�{t�M���¬����%{ZoP�1��4�؛^��L=Rp?܇ި�a�����.3F�Y;!�?�v��(_�|��P�4'�L�K�k�'|���DJ�D�8�A
^<�8���6��+��=A�P�6�^���:�C��L�V�W���bg=����*��IYTT4��]C�%My)
X�m0V�6���}1<хN��"G���>�e�KdG���q��	Z��n���Ś:Y�&wv��q�ޤ@cF��T��30$��?\�� ��Դ4�Ք�X��Qh9I��'��S��hbE�̣#�1+M�L�I�����Kh�<�O��WZ��6;vf�kGS%��̧�fx�|LdLM0�M}���MOb���*�T�����~4*�$�WN��.t�,�w��*��|DU�+�,�c�bm��]�?ŭ�S|7�2�!�����$_�u��sh,}�G� ��E��m����XQ�h�+4��`��	��L˚]1?��L�KfiN��o�.O&_�ϯ���˅���]�s��3]�x���zV\|�c���h�����������"���'yVz��LPwvQ��!D��E'G��3DKK�����I��8�x���q�w2�t���k�6��Z�t���䃊X:��oI�N�դ���6�6�E
�����z<U+��;�Z�n���O�<�"�>i0�BT�h��&��/H̡�d�����(�y�1T)�Τ>��X��ƊOE�?P(��	�*������Ҧ���^X����!��l����Q�l��)�LW&�|��
�l��{=@sw��<Z�;�CF�U-u}d�c�s`.�EKeC ��+:\�,���?޾�' ɘ��v�vۧ�(�PG18ir,������%+����~e3R�6��$䳭t��
��xY[,�g&�8Em)\KRW����u�\�_YZzm�R�_	�h@��:�D���F#Ո�h��k�� "�	��Rb��T�.k�ؒv��% (�܏5(Q;�//d�e�Ak���� Uh�f��T)}���'�Li�@ׄ)B��M�iv�"�K���Ҕ�a5mnp��`��T���k��	8�~������o�~�pT��v��uP������;Lw�����H�Ly!Z�����s�*��V����c�X�p�A~����OQ�c�-��Fj��O_��4�@
�3uEf�1�L�6e<���\)���zf���ǥX;ӟ�ԡγ���ؚ9?j�?H�������L����
e�D�lnU�b��}rM���`�e!�Kp�P*�].�d�!��零�\�N���r
��;|�VH<�̂2;�f}\�1�r*a1%���T��mC����6(�-})R�U��9d�dh�4�$T� ������UA1Kv��&e�5Li�M��-���KM��hkf�~��V��I�0����6��g;wy�/p��ݕ{>�إK��%L��U�7��Z���p͸	K/ncZ<J���ه�9W��Y��NR�哓�\Q��7��5F���qV���sQ�u�=8TQ6PppJ�-�2�oi/}�ͷ��:r ��]�:������k@�w�~V������+qU=ptS�
��=M����q@��*�m��N=M_e�(晣�����;�چ�ܰ�u�{�|�y���K7U���'�0|\�@�~D�+�\,j�� ꫜK�ȟ) ���eyV��m�箕�$v�5Y�L$��P^ _O��>J;m$=k��J�ޜ}(��$L�� [\�7�G��̀s5�!��]�x����-���l�� �I{�E���+��{�T0iyWP:��#��k�͘��0
.�C~�Wy		��n�8]�Ho��y
�(�_�N�����@]ωQZ=����4�L� iT �Ѡ��r�-+Y�,�f{�����&��S�|�&�Ǝ��x(Z2>��d �LrU�^x�5�-�$ lGd�ג����p��^�$a��Vڐ'Tj����0}խ�p���c5�}ě͚J�xY�L�.��@�ic���ӡ6�����"��sW����F��o�P���� ?̇2"ʷ��P���&�M-��i�������T��Gs�����~ڎ=dL���4Ǹ��fC{�]YN2o��<�V�t��͕Zs�9#k�5���Mx�2 R;o��bNj���f�A�TPR���«�٩�8�L<ڱs�AhZ�N�d������;�=�kw�e�A��R���'V��q"W"��b���H�ӻ�3��T��>�SJ��Q��	�mD	�9}:����Y��U �H���O��8d�_��3-nb!:����~(�fI�3ֿ�#������w��t��魗���dl��{F3��3-��.��~wl͊ <���,���'����Zs ���MHO1̴��ny�6�՝���G�8�P�mhf��+�����%/_�+�oHȚ�٣���Y�jP��8�������y�2�b������D\>�C��/�
�����6�����kE>����W���6�Q�������)�}�K��5�!�RZ�y�EV�@_7��pJ|����zKm�u�����J���<�x�@@���=�E.�}S��	�)H�kYroc��X�J�Q�t`qk�68I�%� ��	�r�u���n�A���N��,'Y{}��M�xR/���q�K�>��r����׉'�A��g�mEN����;�9b�1���s��΋�;�0ר���^�]��'�%� .�|��R<�f~�N��%�f[�q����z��k�ԚT�RdW���D�U�����l\1/j$���A��WZ��Ց<�^y>����0>^<�Ħ7Ҙ���E�o�g�B��ӻ<�	p�~.k��]^�v�?{�69]��\�9$ta:V��h(�!wYN����5h�+��@v��O���,�z����D[�mc}�j���՚*Apc�}p�} �.)E�7ʾ�L��3/��+(��(Nk�_T�9��>Ia*���T�����FI����)+(;�A�zoլ!�y�`�8DS-j!N�n����׌� �=��%�P�+��2�3s�.���9�qs_�AOE7)}�jڼ5�@u�8i>��|��ts�r��X��AX|�����J��2*��k^jMRs��Z�+�w=8#[v閦� �a��������ɵf��EHyi���av5Qj�<��w��4�����yǻP�.�-�Q�X���0(4ǈ�"Z{�i�zك�Ӕ�/�1���I`fR�.�r������D!kkբ��;���V�|��[>��"pg2<f��'Ȇ�!�W�I46m��b�(�eA�{ó�]�3jxH֍O������Y���70 /�n�-C�_�&j�l��o��:v�&l"�3��{,-l���!�X�"���{���+��'��&d ��[�w)�ʳ��/.�ߘ͑� �0����^�
o�F_�F�8R֚n��]���|V���΅o�
k>�x�OBX]'��� �����&N�pS*D���x*�]�a2��~Xg�¢T.�Ȟ�C�"��Z�;���k7��>���s�Oa,��W Bh�۫ �J�����XN��6C�W���r,؎@)K0���iŽ��7jU�ʎ���)�c5	��'4K�T�#�#����NFlk�����)�	����� �`j��ǩ��Q�&�9�I;
iʽ�[��e�d��n �����s1h��. ��臭��R��Q��7�LE��#׳�DAF����V�l�ɳ{����<�P]��N�ؼ�&���z�Ft�z�;1��7w�!?��uY���OM�)Q1i�aB���v4��w��;D�gZ����g����X��݄�ja<J���ՙ%���v�����0��t˥��1���J��E�� 8�����(d�0��|�f)C�h�kANzp�����bF��#���R="$�sJn=���B�(8K`/��;�|8]��k�W�c�g�5?,�	E]��h�ա�-�������'p�jAZ���ݛ� ?|��T�B 0�=�1�L�oe��<����i�w�Ȑ�	s,��x��n�.d���+4���� �I�@C�r]e���N*1;��q3��bt���!xN�u��Z���l�$��^U�!Q}���7���M����{Z^^ #Ԍqo�Y���b��Nc�@E��\�8|J�|[܃5L�u���|�9����T>E�*"��K�ȘA�|gQ��
y�h;;m
	�1�(ϻM�E1��E��S�ە��tҤ���G�����n\t��<)#�>FKzZ�����)�2~ʽ1��/c�E@,����#oq�����7�d[T�
FT}�*��Oa���:W��-�G�>�gct�a�w���G+�p'�4UU<,	�T�%B�Y��!`���nr��-�dh�<�g!&��	�h�z�%����GPE�ID�?QKl����Gr�dٌ�P��xh��G���Oȼ�nP制mnA1��/:ܗ��F�R�5:��%\.��7���b�ۧG��^Q��Aj��q%J#��fkv�e-Zm��z_��8<ǌ����	^���?���A�1��$a͋�_�v��ী ��f��t�seZ�Ї�uiMC�_X3_�5?�Q��o
�֖iM�N�|r���8B�ؿ��m� ��f%��h��Pk��P�����{��Tx⤆:>��!|�6ْϔ.�\0��雌���p�ڏZ<���]�N�x�!���HU��1���z�eT7�b�} ��C,��TA<�O�U�{P��K0^R� W!.���8�r�Yj>q�d��a!�U[��nӭVM����xD�z�ԽGeUތ������GW�ʽr�V��/S��I,�'pJ�hc���t�K�#�`�@^�0 :#g{I��*6���^5oI�ŤH݀���(��i	��"������� ŋS�6΀Y�z!*�VEc���/�ɫ������-��6˓d~Rd�i��A�/L\���3�k���8[m�˿��[钍��8
4#�����e�	R��<ýk6H(��#a�f���Q�b���Ǿp���m�a�����0�0�n������&IΖ�ڰ�l�/�ap�R ��p�b9��vv�X�ɝ�O�K��>�\���(M���:a�Sj�e	����q�׹����o��t��Ӱ�����IE?L��	�4���h��u�A,�w)4�5�Ɂ�,��K�p��ȟc����~��W�Ҫ��1\3�A ��U�5�O��p2gY�z��]��3�>�ƒʵ���~�?M��S�l�;G�1���1�Z�y��;�Z��eGIr)�����pU�z��.�l�������G6�w|�q���8䭚��nA ���$�ܖ�����KP��P7�o'�\O{���c�C3�=�u��`�~�xq�5�-��s#�
���P�}�XR���h�ɒ����G�A˭����<���!<��IaG����i*�M��$Ĵ>��SB؛I:۳�W^�u���ZX5�}�L�L�]�U9$���H�S�kE�(Җ��Zw�c�G�����`A��H��!�0�_����Un]y�W��M<����g'�]�ŔR���%����0l�2�S,��߄N�^ӳ�"+�
��x��ť�"���U�����'��v��|�jrT��f��|O�+�{3h&�8��BIMY�'���N�F��(;���'�����B��8�<A�}���6�\NT�>�j^Gb{B��a"^f��qo?�8��a�,����>�sig4����tC� D{o��71�!̇�A-����t�K����(�C-�Cc���!tQ��&_/TFl�(~c��l�>Ԉ](���0��(�a��+Hx	���;����] �Z?�i�̬�@�Y���3��C��Y�%�l*�w��î���51�����Q��y����q8'R0�9��Գ~�+)%�T�#ļ9M�̑���&�>*Scm@F5��h�%`A(�F��l�4�vf`�j��M�;���7P_���$��QG0�m� ;���f���T��_˃�[����}U��z�a��"�X�4_/�6�x���T;��6�g���?v�v��)�{G��'��`8���Pd����ե��g��q'ЉX�+����!FkVy���_�g��<�����s�9_C�!fq�H@��7����6[Hj�:���aI��L�p���G�O~���v��{�u`?#ְ9��r�)�|�"@1�Ӷ?��P�p�Ҵ�3���r�>I�u�k۳����9&��zl鐙�l�H��0������Ć��T�9zb���W�\4�$�Pi��;Aa���u���ZiN����oen<�0�rG)�^BMxA�o���C_�,h��S�l��s��شܠ��}��=�\�ډ琑��Nl?�gu 6�ƯGg�]}t�V6������v�ݩ#h�1[��c��c���٧�R�Æ=h� �k �Uݦ6S;~�^��o1�"8D���u5�����ǌ��Z������ۺ�!�\��O�5�՚.K�/�y��A��5�[���~�ɑ4�I�}�;s�C)�;od+'�f����<>�Y��WX����.�=8��! H.�?D�l#FZ��N��1���=�ϲ��h�c�<ݝ2ՠ�I2�{�9kj �(����F��Ci��v.R��e���*�
jn���z�Ʈ�d~/L
�-W���l��l.l5F�&\�o����/�lΚ�^�wM=�x��u���O��0��V
�om��	 b�!�=t��N��$r]?��u��&��_�&�U���~A�ԑ��M��n%�VQ� +�7�$y���:@����n���X���~�����9|�W��;RRZ��>��Crݫ)>&[�
Vy$��3/��s�'��Lds��	}L�t��}����C�����8�r���3��h	����掑�6ݧ*;E���Tĕ4���);�C�hdm�D_*���xW�1�W�����u3B����:��K���V�Fkf�	H�������)$ؼ#w�1�R�bUO>�
�|]�\�o�U�h�Jh��q0����Pâ��O�����H���(���1�9%�� �%ۢ	x}(#L٨Ѐ�߁�M�,:e���8^�P`ݢz�˙P�.S5r���D����6g�IE��$�
Y7�.żo�,,�ۙ/�E�U�,��}:�����������I�1�(����)�[z�<V&�g��F��1T�V���О
�.��E��7�߈�5$P|�7�L$ �6�,'N��v��^�Hx�Ъ�J�]�Ϋ���.H�
4^���LxlDd��c��+>�Cfٔ�N
���:����J��K�95Y�`�)���]̆�nM�9("�O��b��ͻ�7AVl��Qf�r� ������9��d�0�W$VϚ'-sf��l���f�����DȻ{hɎ�[:^��-�[|�y������s�dw]"I���$���``y��÷Nm����'���8v������~؞�K�Q��ǽU�<5;��޸i\�N6Yk���|4������ϝ��l�ȶ֟(�Q�n��,b����l��'ĘO�#�~��ih�a�TvČ�\L0�s�3B�A����B���I�g\�:���2���� ��}iv�mMjU�f�/�}�sb�9طzm-�ͺ�|�N��҄O�T(� I��Q���9����-2Ơ�5f�2���h��54�TS������W28h4�� 6
�2Z�XZ��N>��������f��7#�-��:��1��V9��^$)5e�E���f��E�.�U�.*,����\�,�Х{�ji+յWۡy(�O����c(���%�\/���)9��}�ȕxx��<˰��c��YU����=�2�P-Q��U�-K�:+*)�(�P�b��Ba�M4v�`_�C������Er�R�r8+s�㰝����'=�Jo�7��y�ϊf"ۯ�f%G7�'K�Ŧ):�Ha.�
M���G,�����T�]���>��H��Y�W��9U��nW0��(E|wX���|	��Ot�W#�`�~j� ԬԬ�' N(�i�P���$9u�XvV�l�>��Y]����/`X�_(DS�>��f�i��I���t4Ƈ�&G�e:W�\Z����$@�'`>6V8m���-�;&�.y�2xI�̴p��H��n�=����d��}�l�8���\CDq�$���K\�ho���&�B�4��W@��)��צ]n�˷q˹k���YI� ������{Ha0�O���<'ptC��0K��Q2�{�[�|��(v:Q�M@Q�w^`H��P�{s^Q~�웇=�Z��c��fZMr��;�<�y��j���Ù�-#D�owzw�og���7&�]G�������v�Uo���lX���d�;�[8�!6n�\5HTgaG/����N���^Ǟj��^>�����˯I��c7�M�9�\�
�*��Ug���9�{�ɹ��i^C�Ŗ|�f�m5z�ҳ���_�y�y�g�œ�V�� y�a�C��_�e Z�q��؟�������La���nHB}���xRt�ZP�c��p�vtӺ ���˞����ɋ{Q������~#1�|�`	"S��@�#+��hb��ԕE�c��H�A�ڂ�@����8Tũ�{�(����-�T�TY�Qo� �����f}~\i-ũh�@���z�G��O�1<�wo�Q�B��э�QQ�2O����g�j����$G����T�љ,4�8na�~ְ�ئ���)c��q�V8c��}��@�ۇ�NQ���X����T�S�mf9���w�ؘZ��C���.�O��`M��3�H9��;h�E	�O����L�"��������mf��ȟNu�(^ؑގt�����Fs5"`�ks.�b�����T���#[}c���{�Ka�J�V�C���x-m?�����U�Ygr��c�Z�!�rN��!���GzQ1,�( �����$݀�6��8��������b_��z�Ѝ*T
�����P)�~̃����niS�ilv���TU�6:�������3ENZ�%z4b��d���F�n��,P�G�B/ثw,NdCφw�:"@����!Q5���P�R�cՁj��^$=
�d��G�[��-!"��*m!��b�ǝ'�=#xWMf�,��L_�,M���Z�m\��f\�������ӌw��o�2O�����~U�D�a4 &�w^�ϒ�����#���|ƽc�\��*n(�G0���֞z����?>wp,��� g�:�NS�C"�I���!�
��_{���J�dP���leY�������2�o}QǕ�����m���^��Ŗ.��p��\��i��;�ʔI����]a��QP%/�����Tޢ�aZ��
�f���Dm�&�}���k~�<��3e�^�[n��Cଁ[Ǜ��JQm��%
���ݔ �)��(�h�K�.�����a��>!7���,sl{���O.��˖E�I�{e̹I*xLΨ��3��`����GU�d� f!�zy@���Of��Xu�{��X*�+l��/ِTY�Q���Keu^�T�L�I#L����$T��cF�f׊ڿ���u*RcnP�[�d��?��Z;=���o?T'�T���U%+(9�c^.˪y�1D�'ɵZ�M8�y���H-��$y�S�C屘�C��n~�=��X��I���Se�Q0�M5�<��l�s�H[����y��������;�ͥ�{`bMT�p�;g^3;F���&�q��ݫ7\1=��Z���=�r�� ��=�&�j�,�����(��0�U,x����_bm��o��D*��ٌ��͓�]�襝��j$�1���s��?�D���L/4�s��`��m�$"�1�u6=iv��Wa^$�lu�Ǫ6��H1vّ"��*���r4J�IQ��9 7Ρ*&�����
fL�jáN�B�SL<�r�RMշBO�royJ�
4�E�J�Be���*���\dR�?��f�֊U�䨬��Ŏ,m奤
x�'���U�lW��A��B�֠D�~4h�Ӑ�n\[�W�Լ'���Ǣk\t�RpC�S�v�E�����L���g�:��c�K�Q�,��~2F�� C��Q��2]/lUs�����PYrE�N����r95�R�읏�kq��"��M2&S3�l��O��N��T���6źP���f��Y��ꪁ{P�
�5'W�? �9��A�ಸ�6�[���1Oۜ�G�x� ��MF�y�U抉�/�ሟ�/�tK�7\Ң3�D��5nM=�,��{Ti`��KK�s]��(��(����n�YT�|�'S)²_Yz\��}X��|�xG���G���3`���.Ǵ�q��r�}�gPx.�<:.ƽj��p�`8�=H����`wѢ�$	/�= �F(�lIE@��-r�OFT{�Ʃ�{�NW3�"�fH�am�#Cl.����Ǫ��欟��\���Y�lry���"�=-I��s�̂�Z{�L�� ��>Y?sO�߻�z"�y(���WC<
W�X�D^U��#��9�0W�Fq��X3K��#M�V��tgNB�m�3��4;��P(:�f���i�6_��4�=m�]Y_��)�(�kP��0��O��+b�)�=�o��CX$��|������K<�X���j��w�1C���毯վcl�s��
��yB4�g`��,��D��R��d~m�.�r1�����}WBP�p�*�h�`=�R�ӎ���\ş8'�}p�K����l>t��*&���mnӥCS�nLj�c|Aa�+�O%3A+�g�*l��U+�1x�@�=���"̲13�"���T0���
J�d�9)�6v���%6R}��h.)r%:��]���x����/�&�SNnl�����FAW��	K���d��`Т2V��Ԙ���m}@��ک�V�ֱ늕�p��_H��01��XU��D!�<��Y4Y����z۵�<\+}��Y-��nG��t����K�,$$������<�f��6l����+>*�Ě�9��Q$l���֡;t_�V��"���=(ɩ�օ���g��:�i�<ui�+`⃘�8���	��Z该��dFvп;��5Sry�i�*(c�Ԕ���E�bmv�מ���p�G4�5� �;�j�D7I|��-�,F���.�I�fNC�]5��R�\J�8�w��Q���A����p��z�3��F����)Z]���cy�� ��#,R]����ln$B��^����k�dl[�����}f+����a�'�6t:�|^���0Q�K�w��L*kY�|ێ��Ū���=a�4 ��_���D+���Ic\cU�P�g?��w[ٌ<[C�C�Y�G�0�V\|&2(BHwbrQ���@N�("k�!"�UC��2����c�������헪I��E/��=q�>�����AH|X��)K�^"�H��^@��t#0ܷ�2F��:��p��WR�W�����މ�ހR~J3�@�m���%� 2�B7\�U���%2d֮�A�-<������� �)h��H�{����j�N�l����u�ł����s[Yރ=�J�'{�Y�����ř�<�d	����/7?�U��1���ʆQ	��r�ՋJ��3�w��S,�5c?K��X�{��ǎ�\�G�	$b'=��E��UG�I�p-s��y��Ծ���2
	��q��Pe�](�A�u�R�B-�z����%�YF�`���d/�v��3�^V)�U�J�.�q��&��fB�޲���Iw\��>�nCBZC��e���?3���B/Pyޢ6W�D�H�[� ��~j����J	2��B�^]�F�٪�SƄ�ڧ�W
0��-�6W�ď�%�{�G�mH�6�G�W_�p�Q�UE�`����#1�6����ؿߴ�uu��i�tv�a0���I*�����c[X��j�)��������#Bs���W6���B�P�f�ɝ�z-�R��w���x��z9.���S�O����\'<r��M�t��;^o>e^�x|��Ye�r�t��\6Y4i�.*~������X'x�|0=�s�6M��?9�����RqKڦ!��%��I� t���Ƌ��o1��)b[�N����W����m��`���?��y��ߎ�f��k>�9�UF�;L�v��-<�
�h�T\�E�欦G�[U����#I˗��,��/#�b�8�_�P�x'�P���ܶ��z��)r�ܟE(`�y�c�D���<��I�{s�d.&u��U`�@J��*V2�ͷF�	�c����l��dn����ڜvHO�a�H���f�<��s.ȃ�&�`Y�?����p޽�/C�����,�Z������΋֫� �`E=Ӎ���H��
��h��V�^�k��<��9���C�%��I���;"qg6N�� �æ�ͩ$��� ��D��A��އ�gy�o�6=�Q���j�_���Q��pO�|�\�ֽ�п&7���L��NE��p�G���]�h�r/xbjR�F ��<���i�4��Vݢ��3=93����>B;���E�M�Epjf����b���frT�Yl���9�$U�ţQ/�2K���4��5�χ���G[ЛG�'��������G�F�֕�1���Q���]�7��G̀�(��c�r�i�٩ӽ�nq���"
�d�pr�Y�.Lʵ�dI�d���?���<b�K���|���M�Z���iG�,���0��,���kqc���6l=���"8�Û,_cN�8�a$cǸ6��n�t���Ϫ;?-<zp�߸8��.�j��4W$l��P}�VL�S�|��j,��g�l�dk������n�a���y��s�)��8[�~�Ҽ#� ���ߵ�\�ya��=3�q�s�MRBN��A�=fKD�\7�dF��أ���W:��F�V��� ��O�";0�d;Y0�R�_� ���"�)�*[?�����VƵ0I�<��&4UNݱ���ħ�%h��ҡ󠫏�jRA��UҷUٿ
8v�A�' <=Y��⽛.W�W��@�����X�sW1���X�g!J08Z��F_b[�f�(2�~���4��b��9�`���p��T���%����6_WXŝ�KI.6���W�H�t!�_
�7~t�^�����Ҡ@)Q�\b��Q�>���x��R*6�y�;�}�T����qQ�1�R������X�d�����5RT�1a�����o;Ija����Զ�Po���,���j-)�+cH-ʟ�K�1�$���*D.��;}?�ZM7����w��lk��3�,��#_�D���9S���/s�/^��>Q8��oX���40�Ӂ�;��(m!x��	I
���X�aS�No>4�R `f+�Q����Q���(���6�'��t�r��<�r�#��$��]��{��: �=�{����o!����� nMh����f����t߲͡|x�"�2
�B���fԄ�����P��YQ�?T3�kp�!D/��!��d�T��ei�q�ʻ�vŃ7���(�S�P�����.Q����JtJ ���[�2	��@��&��}j�X鏔�}�mH�B�C1tŗ����E�!������l��Q�K�!���J���l�RH��:kUgB�#���<�f����us4��>�$/��oH�A�2���ʎk̢�: ^��Th-��g�b;N +�����Y�ʁ��vRs�|�4sV�螘_a�!5/:w�H�jO+��C#���8��<޶L��$}����=�,�'�z��1n2j(|�GM�+��`>*�5���Ib��&#�]%�J5�zj@e�'n�Ҳ���
p����v6�H���vIv�H�/�>M�� �/p3`R���KN�T��Z6�5i@!��������Wd��,�l��f���M�������X��`����M���X!lHCZr˷���(�'SL�$:3�kUIx��Ռ�Jk�g���s>9Hh���,V)E�:ܭ������h���]��ӛmhI���� �NM�y�ei�Q�~ꤴw����F��?���l���4A�:��CN+���Wf^����T8glhRRK�F��9�7�,ѕ��*�"�k��xb�Y3�_��×�ؙD��~؎w��-Y���W�S�ɵ���e��k�+	�:��8��#��ҏt ӯ ���I�2%�f�MJ�b'����>L�T�LZy�3:�Z\^u0�%��U��0���A��[��R��4u�˩5���� �4,�z�h܄����WH�>r�Vܰd��,�#a�A@Z�#�C����d� <�V[?���f4CO=B,;7���	��P����DqO,��
��d�)r�;�Z�F��Y�Kb�2R��Qg��08�w���Q�*ez$r�I����׶i�o�#�iU�ӴAה�ZB*�B�HY��o&(��ӹň�]>�|C�"�"�h3s�,�i*�;��&�[e�rU��F��;�9d�Ca��I�A���P�q5�⽴e�U�R��U�X��Q3���iСK��v xV؞��9Ԃ&m�۴y�txF��V����Zʊa4��T�@���^��3�P������.(�ƅf����R�05����n�x�,Fğ^��<	9	i��I���R��a=#�����!V��x�� 7�x��j�X���ᴯUp+�>�-IW>��(p��#v�B������a���r����S�\���P2�2�ZI�1X���#>?	�^��c�;�`�E�hWQ��Ti��-�C!�t�4�l)�*���i��!t�7e�ܨ\�Q��ϱ�~oc�:]�-���RjD�2�!�����CR-���	���J�q��� ,en���t�y�u��* \��q>�F��tG��+h�A�5�[�!��cf��ʪb0�v�'@F]���?Mj�{8�c �b�m���%��2 3�mrx:�p��G�YI���U6|#�Tm��b?��7�X{��8M��/���=�p��ף'p穵�Gr�_�`s?�<L�.8쇟+�����5�/���%��-���C=���s����p�d8ث�Kp4�g,�R�߻Ub��	